`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dVsprH5u8yMPumln2Y5DOMzoS9kJu2B+zR/ZNhc2AQLY4gLZGJWiY1PQptB+ivO0
00/ZI6S6DpGGL3XCsrf5zCvTNCscAO3OWa8GrfjeOfX6GoxPqiowuI08DRZZLqLB
jt4BRmhKu6YnyV5snp344ykYXp6uGxJFd/4WNjqpEgkcm32ACjoVtXC3tHAiXxiy
RBsVk+Ko/zUjzIwi5li32LcmKYQQo0O9rDQg6q2apV/xciiG5GAsA92lPZRG3c05
msuv7UydrZodgl9gs3zxPdanLOOGIUAkCZ3qjXLEC2B8HkMOZDiI0vB2EjPujM9F
bo0prIW96UiQI5skVKHmlibUTxL7l7o7GxWTW8XbYxejuv1MJ6kp+/ihWE3q5wPy
Ye0TnOrKjgm2nTwb3KBcqMFhqtWn58lAe8C5YQMg4i0MXol/hHuWzLaNwIzSEIHm
JrgM34RUWvv4FOVRS7i81h6iXsNdzmHPD9JVBU4Q2OTKqej8vM/02ps1q2/SPEs2
9HMbkuAmz+UXs5lLQg0JhK9h/fRfAMaBAy2RR9jG7DqaW3kBg3ojmpJUMgmvgyWm
NQJduSP7wdL6NTaUsPsrIVb9NzywFuD4YK7r9Mu6DDPay8h9bgT+eaAHr+Oc4g+A
QrkOp4eOb5hexCKz0JH4ShRF1dxhoIDfPgxcURJlVmJU+PiADfhgbVMRz9vdvUpK
85aldJ3Ndp8hTo6LvwAhCam/QkCuPMdQtugsAeenGE4N4I4gjiu33g11aWsNHeJY
nFd1ipy4EkMMHoAUaASv00SzRbayDOdebfetNZ3fKGeI/SweOhbbv4+BxqG3To15
kMrMza10ivNljkF9HUVXCRtbnPvlYYQ1mbp9mI7UKNqaVw+sIlNke1Ihj5XcVNsz
GHrR6U9QqeQu/EIfhg1WBPOW8dwv0qrN8dIAtoDcNFmSq62/nody0xT9d3aI8hOP
mgbHTay5pFsd98r/PJRyqiay1x4fArKV9CZ2qb3SZj5EVOyCDs8G83Sf8qMfr+Ef
KRV5jEykQYg5Zrx6eLC6SANvAy+g7pPe3SDyaVt64chBtBeuAohnhKRC7TLnvIbR
rHwpmKtMgP+O7Zd88edgSYiU2ly/d5HMN987cTlanxIwcpKMS6sL2bCq3y/so4ev
q2QdW9KaeI0DB9e66bZfhKn8d0FPJpex3uzTxJEA4RwvV7yARL8Y2RmrhNVEMZrK
JqVU8cqoNKeCM6iDUFXPvrKhdjO4N80nY5sMtKJobPGnV6yiYUa7Zq6dK85tYQk3
JZlqYuE/XMr71sBZH/RI6jBB0iqad7ZQ8z97ZLxW2M7QR/x4QXBoWm/GPcx+MhX3
lzk2P7aLg2uwsblQvByQphUuP9qMiXsp/XdmSNtoFfFcQ/oB34dZItF1H+U1suHP
HFjSHqQuQcT25sUYx7zkzx3pFEKnyw+sQykn9ivxijZqqbpEBl8gOZVprjNjoNEz
9p7r21EXePHZJPx+r4kLvPFhye9SQdpOo+lkLZ1bRLVMyKpPT83VezXHnus+QWnM
Hutu6wcR7T0/wlmYnsAIr+Y0oevbsmumgNIGc0TuAnpKkbP7XRe6hKjvJ0+JwNTz
5UhPJy8bgpAxi4xuFnFtyQTu7asUhaOXlRbUWnSTYEHKghv9wqXZGeGbkY0gUkD5
ixPYb4xU6aAw940P0muuHObXM2ZQSq1egAOX6+C5GGAx95VeAgvJ0ePZiQtQ2qrS
2FNmU1M+OdkR0JviLijCgdRKvONY3C+6GVnA/q6Mf28X8VPS7zX6CDuXESCc7WS/
fGZckrSqEwD1rYdMO412E1Ayir4brNyyX8Ia2wuOySYdu5COpLXwd8ltrJqp3XbB
uHL6ZgHd5H5k1mwNagvHlOF8nEotLf9V51HlFSRrzbneGfp1GJMHl+5KmE4C0Qty
TFEn1w4LEq5yUXQKyqKYKL2lgUaqsY3+veiCKS2SGZQbE9C72yxmb8IvD9cixXsL
S3FgGt2NjQJRIOCLmQlNrqebNSjMDsoDfH8/VOpHKC7ztHHSvz/8uY/Ae8ImsHpi
PsL0gxvHJnruSdR0BydxFce3opJewrefnw/8vlO9805v04VmL9EwyrYTvnz9vvsy
6ESdUSCMmW10OQq/RLeUUX31w2J1xP6QWdoKF420sL2gWzxSQEr2m8DHtkffcbnj
zoBoHtTOtxyer/HVSAtoDNuQLclfO+2ZS0aep65a/laOqc6DJKw8YPepcLN0CDUg
R7JfOFBtF3MnEEux0IU9vA==
`protect END_PROTECTED
