`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XYizgxoDrusol0ThKwQnLXZ70t4ieC3Rz6c8JrYMeY5+z5QXqO6VkeftEcmZrad5
ninLaCtxeEzfnvsdAD1fzSYbNzJ2Q6+jc2xFi4JnDpG1CR7v7/CU8qrtHlm61EkX
waZn/RvHbL32b/Al+c0hCZfPak8fze2/9LvfgbeRfrvzxcjVDXCiR/KyLr5l6tTt
nXLnqPB/Wvn7eoQtLVJApf+H8azzxwlZtYlHPd0Tcy7SLcy+DD9kktiGCFFCNn9+
66r2etxKpGeqaoo2v8YJBfvuCLjtpjtFwspHP7CwLFoVq54qWzXq2OoiaGBzQ5te
VNSigMiOQeMSV2+JOLc1JD2NikTh+DqivkHryBnL0D4As3ziZlw/jrJ+AAIzHdaY
Kh+R1XotyLEBomT+1ako9rF9Am7WBPZ3GzQcoNc3Cic83mCvpt5i57I/Pe08TEs6
5tR33op576OekKkivlHgYha2o0QHkIuyQfJeBC0BkxRNGm0cNV8pl3nNOFhtWqxZ
3idxzDJcbCx04CpW9OP0R5ve5x+y+TqcprnDBQBKV24S1I5fhS/wUGuxg54ZTw4W
3UMqHIBvhnU7oGzCg7bzJ/uqC/piy2eSBl6vpAhAt3pJsxkHpl8Mj7Qod9PNnKVZ
TjaiMYT9sIrYO62QmVYnODa6KCdBXsDBN59zKVrsOK/ok/n4cfTy6i05awxpPHr7
Si9sPbz9Jzz4x11YIRHKSVptt2fh96KQiInxQwGof1zSzDht8RVfoYUnjvcSf54w
b4pOfIPVluR8r25xEKU/lVwchb322CBEQGsvvA3KOY/yetxK/LAvD6dBDLHWUFmy
hVAlaDWRUTlOWInD3stBdeLCuEnurw/xlSLwZCxEi7wkoQqKnnik2unIPif1f2Y/
ty3vVeWaH/3TwdHVYRQC4wF2k0wu7WfYaL233Q13NedTuWZwDg5OUdnvQaq8qNme
UPCMEixeqQn0eq0DSwtPeDicOD1AOk74hKbcK+/n3V2fq0jLztJLMtTOVVQc1GEu
Y88OTjXed2P/4qvdhdC1O3ATuBxrXfyH5RN8cv+IV/zmyO86r9sMKO6/8+dwl/J5
FUJdaQ400AXJzQ41nqMFDkS01boEUKikxvKCWGFrgCTsHozU1xye3qfimsBW1E0f
S4vjByDa2BPV+f8r+vjrZXjFoXRDYlNq5rC/2uaYeZxKCpoaVDZe2Vbf6rlIKxzR
2v3VQomvyw9BppYevjUmZ+Wer++YOrT/htPUQHobj71wSb09vn9uGsd7zgKcC9Pp
rtOQG0zCWnc28eqdvP6KW8JdgST/qdgiCF0Zkgrtbo0UwneKDFKNkp2nP3Wp0Pw4
z+IxMz5NcTIRI+YzwwAS0dmzzITZvD6KAfsU7apzSkj25YV3HViq3unynHuTnMsH
xAXwmYtl37HC+8newINj0cwBVPnsASegJYiN0+TQ1odWsRkrOHcGZCTMLce82u1f
2bnVhGvSR951cXnCOt+R5w1eLuwZ+3dikP32LxZTLsCKDVI5Ujllc7Xt00ObTv25
5UxrBNkjVbs1SkX4785yB1yO8qAGbu82kRbIrI+7S4BQco5zpCJXxtGg2pnL0BUf
0OnN5rQ5urs8wx8bVyf4YlDlIqVjFWwuyLn1cSelCdCtMcDKf1gGwkkdcSLEMHM3
xUctYnChA77BQ+lTKCjOLaUWFxZRu3KPlOBmPv5qt5kq/uFJ1eZ7Oii7O9W8aD+y
TQMOsEudcZYinm7G9dsQaUgKZVPP/3KvfKg0LpuA6O/dZHMs+sAiqePW2uGcOD6h
lTEh6eE7/8NV+GT3FFJ4PAy+NuU7ftXOgB00FBMTxhLvKgExIvsOvtdT43jDEJIa
nN03IZ9GL3GnWVE9ZXzE7PQzGTXjEDvllTrFDcqo3M+McamVrSNNNdv6X8APx90q
3AnVlYLBrCRXYike3USKBUdxJ1TRp+fUYN3fmH0jV/sOkOplg8tSFr7uBNeytBMd
FovuZNs86MBDRJsGUJYJssLXcNgnVaNqARIX7smQua944EUDrNw2fFRVqHIz+DJS
vZkaun3ND+HwHB+QyqsKVB6sDs/UGC1uDXGBHsMZE3jXv0ylmO9EpcYN1TPI7Mzo
WC+Q869qOmobTuWOVamE5KYME0lRgpPPEdgFRgCPknbsbTCCkbEfwBIXqBTNhyhk
KnlOTOzqrlXmDEbHTDXydsiseQJzwQ+feJXxCELzHfGye5FHFXtOGKj9yjC3O8Us
tqd169MBElBbsvosmfmC1HvRL03+6Nla50ficrJZkEdekHk0Wifv3FwjTg3Y0eMj
hfilgQYt4hdeZghc0Ml3WA1Ak4Os0z+xEVWPoGSPa7YiKbEEp7r+NSO3GOw8eY6I
IKBTh2dkpMf6ngnV8WIhUhNIE/uyUTY1QmPUi03htmzjd2QAXWh1C08azvcJs8GD
Nn756kFoS8VA2kQl55IkYUug0fi78bkimxPcnBOysk8OBsjVioHvKO5fX4YCGLpb
IH53uRD7n2gWazT5Hm6OMTmqkkWAZBRDEPJLjlz8MdegmtGVLP9Z+MLmQ14aPIhh
STWWpf/d0QuZiGomuTCXbIqNV0tl9YRWe0FxzGDdWkQpK6s6fha8JHjMAEVAC2y1
CczgKU6nDSqfCHqd2GK1j5t57HUB38VJLCikQ/xAGEwESppe0zStFJivE9A7EBNZ
SMc02PgjHoNuA+YR6Y8T7X1O0b5SXDoa2Tf7TNoGF/6CpX1vTlhCv6+NBzS5X8vk
gidr4gO4uVjL8FsGZw27gPYdKFXOH+xiGTo3lDAdG0MSKWB+YBDzZ46RHUQJx/zm
atdKYWZ1e5Tu8zEnlAXe2dP6A7Y060PNNwUt1IFEhHQFavGi3nmdO7FsJ07KdbCX
h8eF2oRIO4HGufqKAC1ZBP3DRtOD7yJ9esmyRw+cpwdESSPXXTSSyUNbp4Px5IXL
axHl5uDo+/rFaPr/GMaUSOtqw+UKX3dLEpBunR/kS2n40q0FktDu9jPzNUwktjO0
H3JZqwYaaHLTfyqfhu54dk5bShWFPFyj+9kzkoeZKZEIIuLCystteBkw7tsonof6
4q5j+NwZeB0F8U8QRdWwN3gl2xW4Pth4ETbre8JrxEr5K/f00La7SREBPyczm4VE
5Qy/o2HHmk2NL+UXc4iSrxtSlHHq3e51WLt42bolnvp70NbcosWSlxhZmKjpQbrl
09apBg4VteQfmMfri6OVdKXnjNP9WTjqMNBg05ADGd3m4eWi2d0x2o8vjOaSYCs5
9jYW9tp/l5p7CaYYNhKPBljAkRGNBWGqdyshbaCcmYgVTEWM1Uy4Hz3+ChP4kT3D
kVh9lE/Q2lIXzjXZaCocMeFYAqOB5YJZ6CykZnIHeOYQ1FmMYGvzIBwo/YNlUq36
ftcW0M1b7E8Zt1psDa8U+Iu8YmagGuYNuoTOqxan5rTez5rBgH+WTqXtUnk+GBTI
/J53ef6ycGtbcJ5UM3f7g4gSHE3KhSefaOuRrCoq/Q/6NLMAOPSiryI+5CRCUv0Q
8zmjwzVIOlvRhThujj2CAwvhkC5STlhdZ6BTH9pCHkhxDWDRjOZq1BPbw8k810sK
O89KL7UIdrgI9O+bfiJ9lruGFuBGFBus/L9Vr4n9uJDEqg/5A1XQZnPGxUDhLI4m
pjf+cUgFOKHEmkeR/h+UJm2wPWiXkqgqyqzRTwwQfV4TAcFZGa/v+g5uQXjGmRrC
8oXYxwGizsQyxRBQI2XAK9nIPxosQc7QpIPLE961NHxG1nwRNpi0YMEQCqGtbqT7
ipGy++e5ln0gqXTKTDGzUHIFUW2L/sVKxZvZfYiGUwPE23WRLf7ZbZtO6os0XkLx
EVLjWMbLu0LQk8YA/Hd+fuH1fIfU3uHquh7q8HUH3yuO0fpj1SYaaNcK5T8PicOm
Ts7k1EQNqpD0h/3vn43sMN3FdWh/q5tXYOCtHACnlAueVEwlqR4to51iD18q7Pfj
aOiZSmpPWw9QjY8KVNUtvozZpp0qiKjH+9NvqfJkbKJLkD9zinp0IiXviWdnBJJW
nJG8XJ0yNZm1MZlwHAuq4KWbjwWezde8GHvzXHOyYtm3XivlrFKUaCXZ4ilSqjLb
kP+c7mE07OV6qZ1JlzmL1oz0ZS/FslHt1AyL9Vm5WecIuKd7LVX1tCCPZdD3UeOZ
oFsAIqNYtoT0TeB4oWGJ09/T/tKzCZkzw51WnKMe3wdZHlVHSFe5OhgDWx9NX5vn
rZhIZrVsulNmb5SU4mEvteLhcgJBdCvl3ZlyUCLjUCQWGjJzDlkWCt5K6ro0r+e9
FonWni8eGiDPIQp6ZW8DAwbDrYMGQ8eS5OMFQ4lXNJf7hwjOwEcUV+5ZWVVeaJhS
x8feozlAH2UA/Na2NRS5ntM3n7VHOATvOBQbXYE1YYVbGDCPUyDpNdtEWl5b3r30
bQ4/M15rFKZF64D/T9pMmsena7c2lXRkTYGoMQ8owLAdkSxQg6bazaALxe/WaJIP
db+r+yGRRJ1qVYdOHJaa0v7yNML+TeH8oYbvv0hjNzhnBX03HCFQMPna8s89ImzL
a6PImjkBISVNsxHNlxkeOL3o8pxkH46diWbYT5YIjkW0rKDFg2yfAVT3mKz5EP8c
KD4JS1BR5kCSqmLudzhTYdn1uYHLCGpFQpyLSggrx+CYyMDFgK3xgClYVQS94J8F
xG0SryWSNZZHJM6VdUvaTEBLpIjbunIBFp7OIb++lrC/puS099W/2EBE8I2eI3CV
zfcDsh0VZ91+51tUYfLZma9+NSYCaFI8eDuEqYlYBXd6r5NvTTwWM/OirRvtl+Uw
jT62ARXL2kEONIi7WEtAp4NsYD9/aYRFCutDdR7q2WszGciiXlCTTeZasilD6QzJ
9bf6t9jhzEzOafmQnr3TnIJ3hCdGDgFiDrUonhCSgUT0r0Jrgbhti09yZJdAiWTL
SKnsvJyAS0iEz4T4IX7M72X012S5cYP7C6Bp4HZnpyKEYzN2YgNd4nNB7mzsHWLj
Vut9ZdLGShvLsmPm2QqQQGrX/yehdOK4Kxc26xjhuqDg+UcTHctB/b2Z3Gf6GOSo
Qte+b8M3Q9fIJO/IDTQ1K5RDj6cbOUah3mI1FXtveeCNgCtABrdCj7pCJg8hhEI+
jA+XWPCmdgdd81KmZO8LFwRy6NTONYBBLjdvwMcJrJyiXt1ny4WxxFgOGWAf8M4o
GVOXBFsY6DDcPVSmZPLlL2tFkHU5M8j32H9h+DKqCvsu6XKafyRmKwMQ2P6klUF1
rfrydZybs3ZIvGCpOsrg3O8W1XryvW9W0bFMHMUAVz2fJ9BLAVOApkmbaWIyg9aA
0XRtKUUK29B/dgTSbPCu7k0FKMsxKOV4ZD7w5QRWgE6jNdrNijaJ8Cvm1mvVPe6+
IHH32LGr0xn/BjFszV7utvRJIJja/MqY7XWtgfIIwu+Eu5CZy0fj3V1OMhvDYvzo
kicW2o92+uYX6+OYG2YRLyHNyDThTL3fEMmn52rtgcb2Rs+5275+81/24PxzIpbF
wvgkRYjxf7nA/6LzWmK2t1hCQdnrcZNCtq6NbCpdD2bCr+HdLdS5FVf4rum0HK92
tKglLlEf5vZhH0wTYCj961uyRjeY+oipOGbCI37FY9xFzEiZDuHvRHuhi+Yp4hz0
biRjwg5aRvZZF3pH7GCp+qJTxUCFfMEDcfbUMP6olDJ2HjP5kvURiOpE4ujenX+e
E9AYwLmTGNPwj+Jtv/iqqGMR8bFzouSG7mNYA9GCVzPI7NfRrqkwYgB1SLHCQN8+
Gtz34FyMFRjOjtxiw9524txVk3sZXdUeg/WtfPX1k2L96NMzDInW293IjlfQl8gX
Aq1uCzoaTu61uTd4O9EosehwJTKTbmuvr2xEjT0Fe+9JeNA7xQ+K5M4GNn672gRW
I3AqdOEMJ0ArGb4hbZmpoYi+uCS/YHr33MQ/xUQ5InZYVOK0xFcLP+8LX6a/N7ym
o4/IMlbCvNBIDbMTLzsDa2pbATkoHbLQaqFQH4DLJ+dJpC6mXnL/ojJPXehnoqSr
jFNgkF0hCecugN/yWuYrv4Lx8t6H7MHJfnzsEn1+z5Q36Uivz06uxnXybXLjpvBH
32lgm0Xn+QpG44bxW/6d1rOlUygdLm60aE1otSbJ3VYc8rw9kcwHQw+zU8EkzL1Y
BkM058UN8LTmpe9bormyBVuFAerhf9K1FzV28b1poAoPVha3nZKh/qgoo6yH+crL
vZfHxExb4xa78sKHH4dVlnMh1GDjfh+G1aafynA1/ticVJfJ70dZSpZd6u3NzEji
/bzQZUQJmq6LwhlWL+dNjP3uia0cZ3hr/mcZaoZPVxjAczvFymnOblPNTse5cDGF
ZABrV2tfV2AaUQ7YJpAyOK/GU6uBKGRihla90V7oyRyCeOOVoklCxpWErnLNixp1
cHnNAHy9VRPJfFuNgVLTh33/hEtg+B1LQPCUa9okb8trsv/4Ufgxu9UmpYZuNLq3
+ipH2iQa3mhm9okn5+G5BezUhA5T3euZScA9rL6qC1lMoCQevCWGgdk8T0IB1TGQ
6Mfq8cOodxxoC+bJpJutd3SZvxiJfhBYGdCboF/w3Yq1xPPUjecOVFHEkF5dBMIW
w5sm9wX1hqMXf6r4hqWpvr+IE8tVHIzcjkVSFCSI7ueUAEKrX+kNGYRwqogONyo3
NcN1GbkoyqvVz5vWwl786XJLsmZa2INRBemeb3S3fdPxaTKSI/cYNl7vig2tHJlI
u/oKY4NzPPCGgycykjvPHJPqeYRRmbs+BfOpXpN31NC6QN91z+M2jVubtMQ1cieO
xYMUXDPu+c+D5+uXbHE5Jbj4h4z2cMiQJoB0ASd7pMQ/Nk69pjaSKxLqimK5AZoh
BCytmvitZ/rXvF00BuZA5pdyRhBQg8O1Oba6+hrP5u6U7mEZaHFMeBXC0ikm+IeV
XBp8etjCQwjEZWVqF9/Ro+GSXvLAVI5Ny0ZdlLjl63SC225oMfG9LKuFwCVWPUls
ZbbMQCul02eakVon7dr6J0Ld1Gt67zyJ7aNfrnuVH1mZ75mV2Bu543vQm2X5xcXh
1hsPVyulKvQylfZw9zjmiGI3h1FFb8rf7/sQcY3xahmg0+GKOcZ2e4aPWwlMNlfW
W4AgTEz7TZQmM+zwjbeUqgzlAVEUv+uFYR0e0mOdMxTuZy9Y8TZFudpsLmxg37dt
aEAjuSkZZRlkfXLPixEBeypo9rxxk3sYWgoIm/QNxzeMShrfDy+XtAS2ZGpbVhhE
vyXRmSzc3qPp9NqCivX01AWAVhSzIuLZbDttshUzqtaUOd+zt3Gv0Wt2OtKTJsrD
myNnFI2pPwrOV47JB6CpKRt33wOVVEZxROORmIv1e8uGEJG489/D9vabXot9EIsa
ZrSpSjPhWR4RwnJtKlVBgnbkvHDPEjf2c+VmxD1azVLoJBYScOvoi35hB6Y/Ut6w
8MASC48RUusaaf69K3YlZpjzm/bHB/s/YS1YR6WIHaXuKrxCX1nLQ2S+DgycLxob
iNdsHgR90QEEUNlcWN4Y9XEl+LJThynP84lHAKzorrbn4/XXmiypjC/UTTvq2Ppf
XLnaaWvLbdAoZmTL/Rvce/PC9mJIUAzpE9tt9qWV2p0PnshAJf+FGPVEIMmCn+8g
j78FuivywidBnmhcfRLwZA4hwHRefDX2bd4WCw9Rs3j4gHSYrU9GImHQvx2nbpm6
m0k8td6Ms0H+dFkdKVMYPUEWhNvn9DNj6o9s3fmtui4difBxRjRMawxvTDfGW1vM
eez4f9aCWeSaWptiXZ3yqNLbbA73BqXm3pNBpaChZ0RYPlsmz9Vc+ZemphjINeBU
//ebXrPjrd8PVvXiAW245IDrlz7iIyggHT1ieUgYymgLiZ/uFUaGwICXZ0kALIjZ
hUikQnvOfnx6S7Slt+zxf3b99QVi/FDZvWNezciydPPsP6BghehNwG8wzQKnlJ3J
Cbc3gv+5HR11X6htvhxHMOM9AZ3u3DhsUdkIuZzbzI9LdOOaucWjcJJfwCX6QTnE
29Bo9dgWSguYM3qKVlc8tujHQdQWkNZbuxD4Qp7RkXdOXfMY3oUI3MbbalH0RUrs
0HXQjEQwORbfJ930Fw2WORKvPwXkGo7jJDArAhl7Zkj0dk6HbI/2z1Xe+RFjxJbc
pkhScLKSdY7fOFX/UW4exJeNi4mnSY/LVAbOWInLDXAZp7qRjqmB5CeNuOY2I6gP
vdvr1+HSSFNvbENq0iIDyFzMFuY5zdeMcIS5aCIW5PyuM+fKo3RBIh6Vae/WQnvx
NbsTHhCAW8x5moR5tRC7foIrgIrbCjCh8qO3qQ6VsfKR7Y4kqot/ACWOtWbonyNE
gUVR+3nY6BYv22frZ9or57TItJ/DjDff5lEslVb7I/eby96wwuj0XSXQSwoo13xZ
NMTCYGsyDafANm5dcJdMdR1cg1EAH9N1lo21gWkwETt+ZvT8gcVzM1iGI4r0L/te
9F8wsLYVJgRk7Vr5cpBtUhEM7urLcgR2jTK1N2u7R2a51vrDbouvu1WZvSzcMjxH
YSqSp29kXW7lS8IHDkXZbtCAFxJ2JurPRLSB+XVEfP+iLY0E89+zkvhh+7kwH1Q1
onQJGxelsV10Q9ocxBYuY9cz4g74b/XdLid0ZuW8Q31nN8qbNbI9T+b5T2rNpnAo
BRoiUwjmp8y5aw2Y8p6I1UM3OZW3dIc9cbC9Bk0HaU72GnXoN9t5TrFWuHQpetTy
vQAJx5xiouhdRuk/Su7l0qA/aqGDpMG+kg5J2okDKMSJTo+jLKIrRiqAThF42c10
W+Z3v3adiQuP8nuA13/hQ61gECUp0C/BNvKX17yRGEeCy53QV6EZN3j1WnoxDGQv
1JSTXPgxVuErniIGf9TUqkdmKupujhMuuisybUJjAq6mTnNCVNj0MQxNbXvtn0dT
lQAXMimzrUFmNBcLy6yiw5AjyUOEJ5B9lkDPn8tKotU=
`protect END_PROTECTED
