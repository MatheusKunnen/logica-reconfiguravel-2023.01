`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
duAWAkwoi61HkE8hmjQFqksuL19TDH/Rvr/F1PJYIPCm6Zptfo2zj82aEzoPKewd
/7dV/dJTOOas0Bu66ZJoBDkvw1JyJibzrEjxmckUUVhij4kunILSeNeCcdJySaz9
ewzkdEF/TmJ/5NmAWHiRkZfPBTYJCpI8C879GIGFd29KZwBgIW65lxGtqmqkppT8
Wy6cPgfLegA/f0uLS1AIlAYkZFfOg9EMrJAx1SFIGvwU4r5HfsZsgp4YV5nKqV/G
JMC6H+hBtqVj1urAYzvXIB/gdxC3OWk6+J+1SoplDsovT8eponmtSnYg+B9VqGp3
WkCdM5tQcHsopbDkfJwF8qIOocwSE9hoWp8GkbrfnXIQBvOUCT946n3+TcOQodWY
fHBH+unuN9OqmS/iod4mJ4nKkf31F7A3nQNThi1rQyx40kIUm09NcbCWSSEArGIR
3PUmokgI6NCz5PdVcGLCRYItAPNuDbvYo28L4O4xgjFzkeRC6KGw35sjKsDQCm04
4XLj2Yzi2NJML3EBhTna3qCDW0EXKTLZ55jBXrSNzNaal+tSvMjH/eT+Ur64siKT
eXavoRXtaRuWAw4y13K7Ea3cBNtEeQ8rYSnICijDMtikw1buQnOqVw6yb9Eg/8ii
7iTr1mKYEeHXhBVgInqJlptVBewfbfGEnqQ3o3cyb9ivimdSuhMbcEiq1rLcZPyZ
`protect END_PROTECTED
