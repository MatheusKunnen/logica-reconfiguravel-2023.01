`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZDnVIT+iaKO9kyffjj8A2Io04pOPTgI0c2HycnCtnghATuKkusHaPblbp/75M/t
Fkb0OuJuvrtnTyMKlIhL6lCzIsQbL/JS2SGs9UZuwspt4KCsTRwTnIwmrzXaOQXS
988mLh1Ej+4bFeMzfjX7dnYnefTmKtVmIXT+geUHJSz6u7Ri8vM23rvbI8ZeBAbN
bFAkt0PPlW5MNLdoNaC2mWyNhxhEFAHy7SYyniOU2RofRR5/ipFPKW7fAIWmrdo5
ud3vLDY8liqqM0XuJst5hRFjkdhu1IxjZP51seuVIgszwJ5YPc45HGnKTcIuPEJl
TC911qPXimaY8EULWrKw6lv5kVCBsZa3yN8IRYlsdjCabvQgOiWLKnTljQ6upOIH
fsvImDySI7GoS1bKBTH2zTm9z8Z1BolnEmHCq2qOfcWUSoJgEE1XlDGJSrwYW4/6
kV+V+6avX33RgJqGTTwbyutKlnWlT8SxgkNm0biorT3eApFe3lxOf7RwNGlXRckh
lZqmppaR8HJmmTJdj29BCsNbklEP7XqypsmFFyGSjzQnv+t0WKODON2QPX0pqodX
ZA15kOYnF3TlyZvP1qmH5qoi9fift/CgpA+vJ3RzrU2Sw2FvcFsZ69ptREoeNINf
Fh8WSRGwW4GLDmNqdm5F0w==
`protect END_PROTECTED
