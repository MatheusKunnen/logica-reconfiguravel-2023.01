`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BoOZmDxrWAJD+2XGgHl4eL3wyrTpJanxFxJb31tak0zoqagRe2dAkG+QIAbdls6h
IehPW4MGpVQfB+XgiTI3ElOmTcGErsjzBNd/xqf0rJRpR26x0XDNOHg+ccNB+OdU
aOLwFtQPEB4BIhiHBpRTJy2C+S+2riMyYdkyOi5K0NpBqUqvwHqRHulVWdd1f8wl
P/L7ZcpyCuKIqpl5HOSgEKSObuRpZ3t3RlUr+rFAYQFa8MXkFAzeFPr0RIg4OZiR
zzxF8CQWf6TaCaHRWBDd7HvytH7+UR9aMZIKdrphR7XKRNquF+GMOSYZb3GsGgL7
S0IU1HgOz+uZQeLtwL2sI5asKzSMA3Sz0pohVg7jShvvp8BoTFLdKjf21fnKJUTI
F94iCJSzqZI6cFPmBHu9HPAHHU6pDsfbkoETX3ENr0j8U8W8YnWNTVnC95hRphWt
IWP5K/hvLf4aGT1YT3I920KG+9OJeQzWkUYCtQzTc9Y3A2AlimzyCGtw23TkuJ30
ll31AoIcLx7qd3M6aNS+jBmiSuIEJL8pPt4Jfm6CDKL91L2GzHzGUKyUgiBoZQ+H
q6Fpro+drDh5aViZnxI+w2Duof9QvdhZi/y5UUbzk+EYgzSA6UBUlR1eRYtzY7v7
4e7JZ9gShuaekbqhTddMz5A0VFUCRCR34XRUZ7dSMxRqWmLNqD4+PsbZu9zMaX5b
v9KMOh/BkIwePgJBUDFL5H+m3IcrHoEy3VG7bMTgvNWzTYTSRmGz2gWFGQ0m/dvS
3R6kkgTYdZK+Uof2r3B0pKcdVGAKZA1R4/yWObM1/LY49SIMqiabG+wNpDonzsoN
qLkc2zgvZS4/2/Ie3TCJ4TGtIctmrDm+UQdwq6FO1dUzIelbIykAsaOOtiJfdNh0
uApogPPydyjqFWmowREKzhDS1amlC8EQqTz63vlC4FwVfmkTpMv2ZNLzGb/nR0yE
ebt2fEnefW5iWhx0mN37sHyhcKoRDK7PrOyHqCF6HRmIvMOb1ERT41YZhFH8wQPA
GDgW6737LVlZrqNjY1vmcnnp2zgpUuO5pVCNk+718jMZ5pTHS2O/oNM0RuihTqqf
FFRzqiDFZ5mZrv+XKrllwvi8HxPbS53NHu8L5RuX3aOvM7CdPGV4ZGV2tVLK/jl9
T/0GgqIoEx43o4xHfuoZfnbtaIy6ggsrTbBPIc/gg8mIKtlj5xHjzEq3ZrEfolLM
5UlypoyoBvKISa24DPzJUm8gla7gHnQb47+NIVBoPtbkbyIRrdrhxi1521diHXnt
ZLhpMhZdp8ylHP9yRC0vSGVPqJpaClG48ij0qpA/8smKD1Rd7GrYcew6KTJNVUCv
Rt70T/0yw3D0mqbBXsXCWXEm2N5reF4GRT6FXfz48gb34GJFMWMRzfojn77LPiCg
EXZZ6zhCvU/AfXEJlRhI6ju2JGHHjcxiUK49D39NynT3JYbK8XDdsRV7FeBDxh+b
06UyJMUEhenUWBdDQ6mL7Ue4Ct33fDhKyocu8UP9XpYamSg2eMcXjlFoKPJvWDAZ
RG8BVJdfhCL1TRURcS3/1yaEkt7VuRZSzE4zbePAb6hacupCNXb+68BmPf7t/eoS
Dv8rF4s3XmTqkycpc9HefN/L+mXlawS8KQOWRKy/g7K+a170lYXGi9U1w9yNlTAk
MvM/VEMptmS792XgB8SvQ33GeuPpC9Ga/ea5PJz+bqhN4TtdaRPtKUP76eQqzey5
42vC0LborsgmNqf814Z4bbcD0iDicAm18Vtgw5mAySniJ2OAaKohTMEhwwpjb2T8
H5E6fSoN4Qrh+0cNynuo3VuGXh63mdiL8wqUwYWr91gS+zKBegZhOh8PcFYkiYun
gUS5fZJdZViYDelqeYngcEnA1aldOihBGi9Lzf7VPNAXFJ6+9XLUMNf92L1dmx5B
9hKeRCBGUvvg079W7PKYX/xGaWN36ZBwYcCEeDHeifq7HagBJbfzLcEQTSiZturY
Uppp4yTEOupL3XmP2PCqZJuwF/4nnOPxJ+SULzA4GRKfvXHhFOOqz0rtDCwh4cGC
ygOe667wuzesdWplN7+MDq518CPfc3/F+rYSn8hqKyu49zxUfNGJHkMgvquyfL95
02JyRP/DWg8PwyFcuSrnPHuQW+Tpy1wzlOId5AM6zh9pvSXMeqwoTPEEeKUGcIxO
7LapPKEIYHkkZxWsy28ieTvkiqsgIyAXoQ801m5olVaHBd9cgIkW2qxZOXae9Qur
rNfk6csE6QaqijNdm9ldIfedGD+dWajk6t9VV+V7MFaHVOrc0WNX2Wgcz5upxPQt
Szj9DWR0i+9SdW9HsA/xHLv7NdiuX7O2sGre+YBvRE1WxTFMDGHHN0vYEWqJ8sM1
Zg++Q2SUn4TuOui7nO8KRVfxJHPlruYytwrf7CkIbvcDQUt5pYoFQwyshjqS3E4/
3YxrpD4bOSb0UT630NvNXqGQbta28P1dVpzfqu3qh6oH8ezCip/SkD17fIGffAWu
sbJyRzqeD97TIGc6qamVYym2R58JR4CDndEwql8qWJyeJnALoLDlN/JPJCquKuii
lmtRXgUJ6ALOE3P511q1d2Ppq2RdcXj3HE7uYN8ovy0itGr8wyXJ2vZ2NPgNeKr7
dgGhYX+3bVNM+JAagPQpo241k0/gejIh7+7Y0sahztOXhytxJAikYOJY3fdTdWHt
n6VU1YP3b8Q/2fMnvJSeedlbF2Ixa7/e/Rp/aO4wMO2Hud8CCnHrgDOfql+GDzPE
mqcN1iXcYJSAoNVvlhBu6UIV6jlJB3j+oYoyjF0dlMct7fT3qe0/DDOg6re+rrTN
MNdCZNejSzHaikdNxzuUpsE8kVtT1GJG/DddbjMWhSIC/oVxi0vNsioWrJOswFBa
zfAY0V5T3frvUX6fCmMUZz5D8r+MupLGQotK6TCjdMfbcVGoYyqy7rbwcubynWS0
UOpoXdDomFf8SK14YjyEK7qcXdDkhQs0dn6oJH30obX2kGB1WStu7KrROcAnLwi3
v6wBgqrFjA56+wT1eknsbWkPGxT9GRA0knsQsL1pqh4l8wqh2M7hkvJ81ClOAGns
WNyrEx715fRPcneov3a8EfiVv2cUCs7BEDY5ssDVehAYASmKjU+YxJ4cVW/OKh93
ycJj4XirI6Z18+dd4OgVndRMZM8SGNove39c+KAFQ4OUqCWQsrFqT8QJBAijBY/+
dTwgGd3+h0Zj6V516ZkmzdOwVCtF7lPzF+17aeRyFg1cAfc19retOvw5mtLx01Id
nZ6b5UdhgVgOGWI1Zsgl/OjIdmzjYMkNNB8vF7FMBfrTx9qM8HKbi+jxiyKelHP2
usMP5tDcll6DEvToj780/k3CcP2lMXu00vxmeHPiWwz7ipjQbXR0Rfv5RA0DHvDu
Ey4X66a3BI5t7PBPezFMSdcOHxBnaCmwyNgcaoyOvuVm55l5iznPZ/B13ymCgFPM
x8hVXf5IJ+s3FB99u0uV87hmqjkcMMJOkdHdqIMS929+3s6kShZ8UZRIUiD5m3xq
FHX5gU/9vjl7BPm6Gpn1CbyMDs26b663hjw4kTJx0UI5wE/J8nZNVxjiQ5CFQbiK
XYdhY/3nKwchk+HbrN32nKbzfUJB48IIu0Rfaf+/jJL9VDeuTS/pEp9S+CU670kO
9vIymGPsOxFpZYYglqgiYSnoQUKRWlbvG6NtTANPmuX4U067/XeTH+UEUrub6L0v
r9JdfEze2MuA4sJWUxpAWGYdeE05tPY/RLPa/x/MF0yOLZF9/uTwQ6cj/j1kDkME
iC0vI/jy3JyYWkKH4hWFKgwYF3DESmzkqOIiL+PoNiD5cPI/cG17w2bdSmBSvAhU
KgDeD2n0mzDxJDLX+RNlWDskP7gwPYL7V+p2mIxZ3Sm/DvtnBFtwL0Lcm6PPtHCi
30o20/e7hphCAe9TJjRAwxYZMtnBJpbeeKC3RH/0P/38PjTvXipRpLrhGdUqCO0J
Civ5PNymllDTDW9jFrFPXqtwCfnB56s5OKUIFTQeBZRMXfaZZyMvk7w6vRwVljmp
A1OjveBtWJKpnn7lo8MKlWC3fXre/1dKDQGF9eFM8/dHLAmJay5+DHAp5eggOarT
aKjV3OUK3410DXqfS9LxGepQkAj49Z7nIHhhuCeti5shpUEMe0rAu+xaIhbaUk2U
wh9nH1NeLkacF26g0fHTnl4iOsuYKQPSVbZeDzHPQe+1CprX+7XKme1XeuJbf0fQ
J9XUjXwQZC6ylPpTAJONW4a7MX9NJZn6XyXDWMtGu/fNQqjL9eg7Jm6HqVhekk9I
Xof/hzyoND6nJZI8mhXxVsjfr5jqdn59F/vAQpQtrrbMWOvwoh2U1R7Xs4h2FFF3
9cNP3wKxUt8MjsAmICu+VRJmLSpbjDoiFNvgsM6zJ5KDCEYzfiEBvY/B9EV1OA2K
nvwIBCV9/OQg+ZJsk80dpu86xXvVKQDryC718NJKjTYsNScWgNq/qf1rv8k0B7n5
3pkX4x3o13Nz6gntvTznj1S0AcrvoG9/hnaIE3jnI56yfvPLV5X0XZc0qzu4wPhe
ufLnkz7FMWDhCv1WtwQdsnxU7Zhs2KZLvUGSs4/Jly7w9UoLpUEY+Tpzn300k5mt
MDVIRoiepF7pPu6ls5Gfh/xYl3pF+7JsOd3Jad/EenGksGnT/3mp/WC57j7gb/rf
9f7qTSCXzfXQP6yfyDmq+fyTwm2l0ukpZpHV4XtuHnYyJc1/x1wq/HU87JwldJWN
+zVIxQrsWsMQiE94wtobAM2XgUflal4a8HMb44z4BvFHEEoYLxKAD4JxNK9Ewjmi
pv/8Xnnc2YqyrhF8kzzwckhomug8OtLC+bq1X9cJftBM5SRRyjCq2sj7CqazOxQ4
qKZnq9wHHA/nI20hpmnUohci4eNf+3hdkDd/rz1SMkCXFsF2QKY0AU4hP2HBUfDD
ndfNrvRLVXLrRGqAFni8zmEJ77kxYzsNHqZEX59YvxvbnAd/+nqdiVqG0EnBAL0D
sCz+T2l3CKdHOdmTrLr6JSXx25x1dk9b5TNl2Y2ecGR0J7lq0tRYCDhGl0FPwqKr
XLHMxegOS7Shfh1TrTN0OhbuQPiXs17+9tpQStvj9iqLzrELe4HJZ+tMDNTIXIzS
C/4seSng11mG8oiayRK14HFKCu6eLPTMbTSVfC/1wXGKD3PDX8eMHx104VrSsmqc
8m7dhMSdfAWgxfuED4bGZfo+PabGP9agC7e2tbk4cO1F/N00EUWAfAX+ZlPOslVl
2m/kboiPOVdgeWkfIeDeyCaulqAAulEUrADu1qI4jtMYjNnLNEQqIK+6LZblWIxp
tDCzMC01YSPjbotoXCEW9Zyhcav01pUAOY88FBorkElS63o75bLxUY1z5+1MGCgY
OpDborf5f+9pDfivDLoUwiSfRUc956B7r3lUQp9+FRSLi2kqSKxUv4qhZJlBGYGZ
pBl5PMitlsRBeP5zVxxNzDbsmd5YHnJpf9V6X+kewHTISMEtn1K3fH+bdzWgHrst
u97t83d8JnneDCKDxFi1Au/+9T13NuNZimwOVemH3YfFpPfLd/KaFwy/nP+naHT/
s0axqpcJIaSx4rTk5+x0CelNiH/Ov6kLawRYojLvLrIF/Q3GX8Fwg64M1TRJywls
syvoKekRjkoY9lingmvBebdtvAb6IbbdtwMKLiBvw7vyTr6prqx58lZjUUAYh9fC
31XntTHvtGzoPZWU1aeF6ZA6qh4JOxcFiSDuD0Xvgqdn7pQA1KSsPQ7ARaYgDzpF
G8pWnWMUrE00MFNZqQGqcTgdLkVdRa3OlX5KgQiK11Ntc02pilBYn9a/ywwptVEz
TePKRJVhjTOuSY8zy6PUGP58rAmNwTVqaSuwHUVOCcupsW95kRjWiSmGHHcl58hu
bSPSBXsPxtmq0Rfndnuh2B7WSxp5udYYVKVP80fW1v2MfWGHV1WAMhH+NwSKYXU7
tSoho6L0Y8MVDBB5DTaJ39ehdCpfEdzMzlkwI8zoyLcxlIkSSz3wXOT+Il25iCiV
9gLRMIkcwpHscLDGrk7HrRL75qNjB08xadf+35mwu7/YmkpPA0hS2YwK90VgFx/E
WsAk7llO7eTfTSO0N7l1B6/bUspzFASqNdCBG2fNZEokzFd06yWMgNnMUwIdDaKD
WtQS6QNmwg9Q3wkKh2FPSuWtZ6pBBm+FmcIwNJpBYlAhxIrtYNqXorIobsS6c50b
VnS3S6xP18UzDQTbwSjSuaZ3eEtTA+0YEJQnFfHmyQj0kaXC9i2HHvOZlr59D/vx
8fvgY9ms0UyeBK8Z5VMw900jV/zDI2WfrdXv3Cc1unJGIxzaLMy7EkYU1C6rm6yC
6hslg57Aih/3fqhIoI/+dnqR/90dNTb/FNulawMjD8pZKLE7gi9mB+7C+UkOBRMv
Gd4p8LyFQacykvZZ/7c58GUBOjWc/JoZyy9d8OyCEztVL1fkpw8flGbwpqtzufv/
iNQRTcBEZVuytXquJbheJegRJXHcTuilFwhucDc1oGwNMkL5LUT0sxxCuAmaodVf
OVpFNWRq/sv4R7Mto4MU3svBd4aOa06foCfZ6FFjbefM16feavHUKRnonOZu33xx
QBMxV8l5YQVvJ9l6r68DAjtIwXJIS3IOVAwMHFwx6O6bzzOb97YrFgfo33/5DkOb
BTA36TX+hq779nU2s0Ah2FnKNeiHBRaHUzaPPBfcXDo+/Ib3q0LFVo2W88H3lTZs
0MNjX1d5RofFvA0XEN0rdkeHnCcxNGPgn1MFGAwKsDkZhK8NWuXi/bkcVkPHSDJd
vQJCjrwJVnpFtkVqCVcHrhbeMacrtK6WkQh+CXatCKuizMeW1neW0ZkfKbThXFeR
QqPTeLGYHKkA0Lt+Pp+jtJcfEtYcubEHS+ZCQo9dSmET6LJuA71HljyWETz9pQQg
ojUUwbGN45tijdatdXHX3SLmS1A+YEMKGm8fpme8xMZZ+bpzZNysuMfLBHxVTyH9
wazkXc2Mf+F1MYwF9yyiMI5qywrdCFQcvARgbMkj/BGtod0PNS6mnsKyAqF+rCDc
afxwZCkNkBI114gCA57kmhCWvXsHbTKcs1lAsYJY/8RyvoVW6cIGZ8sRgwFAmr/i
mO9B/MrZCJrZbu28jyHZSB0DEh5dm6ZKtv0g02B9grYpsitLj5XbO9eHblF1GYpN
HECG7339y0Fd3dCdEcZ0TDQ6yIPsoeuI9vvoOTmT7UCIqP/dsKGi8Fxb03SOMV7S
IdM8b+WbVmMAzkY8iquYl8nTAANJtLmwViEZajs9bvFIoT4ZU+/t284nbYhnFaeB
GRtyix0F5OdqpVbLIrDwuJMFQCKmQQWROkWU+CksxotZArxRwhYDdvrOnQIJwACb
zJo2/l06TDuIt9I/LOP9qDGn7H35xUqcgi7390hnun20r25xlCmh3glyf2FM7yeo
0YxNPj++iNMXZc45S8duW+I6E2kfCc9WwMvUUc6ZJwzB1QwcA+65vqKfAa9Mp24h
gwkdtCkycEotOAT5emFz6xHq8bG0s3r5weEKMzZoJttwv24Uz6WJfKJSI7boKu4i
m3g8AZP3sOrJPLkS5WNTCBZmH9X0B9YCRe+fHl1M4UDtJlS8NaZwnOOZ5jOrkfcT
Ht3Od3h5wUBdApw5m3uINOkHjEw6nmWTCp9lcZbllqyYKiga/fJIVelGprwmoExk
jOxH7kbVH0AoloQr5z6DOtuLhFtKx9AcEmDYIxNIKQUDjMucp8lGg9xY+Fx7U7bC
NERSPcWGFmARDwjrAiUpHSVsh5zoUFjoZNLvwYe2SxXNQbmgwpDv4387mQGbjbay
AtKwCJfPsMswFsgDyWZtCUfcFRUmxjFutoFWb0P2z9oLTH7pC7oslaA0tcM8JmC0
qa+aWF0H9Joxy/Ed/NgTxZyI/ouxt3XvUQAl7ePgZpgC2luGY/ncNseyo6sGAFz+
qgfky3fdVFQrkBGru4jpHooSd+5KWwCH30EsvlXNJRzJl/WyEGOQoBd8F6Zh5zmt
IOevRhK9t+WsDxdqnslsPCf2fPsLkHLwp4CnotWMqcH5Ivp+NXtDxOp5o8QXnpYn
JPDeWNjnMrPsbDbmfiaJZT6pBJDmYB3UIYBDhOod9VrUyt/srQR1EpZyVTnaEXzs
DtDRxPf0nNn2rwXT4+qByJILCRD5sabkLN3ZNQRf1O88nCEZoAp1UK/fWS/RDazC
Cm99tWQmsUV67UypVD32XP8LGFkzDFBnVBQ1SGL1SMvPkPkJ8o7x2OPAmS2dANze
3JdpVvfpJP/r5xuJjGPhiESpdHZrb/NlYVKb+xGFmperDQ1zCxZlnLb+fpmY40un
CeVx0cTJ6viodMuJvwSQ7ArpjENEied6aK+OFJdJwnAlZJxsQTSZPXlSt5oc0o1H
9635lGGsbn0kT/HzIUTa6g2WxUfUWmZhn3KhmDj3EdCXqtdD+jLfp81d5/ZY9sJ8
OTR3ZsUwjO/ySdRimvR+py/k+Qks2t2HxidybJe2366sVWEzxlxYGdzYtnON/+/N
kdlcDwbjsFMwK+gjsr1aWtdCCEKltkxe46ayhw7X4EsSn0Vl3J1J+anSu8ypGlLI
DLOecAB8GIvWcCLSZhsy3n1SisBS4l4e3GgNRt6vhSO2IGSfuI7Mq56Tr/adrHeg
+zG8gNGEUomnuq1YUQdIciKlZq9n+rNHTTEdAkYPlJLC9abnHF9Tk6CNijr6Bs7S
2Qjd7KOvi/hZHZW3B133oIYaoUgLO4AW4fwjKgn+Ly4rM8gqt9gwsaXBAjaL0oEK
kQhPgd5MnVNHprEf9cF+ZBdE4YeWTr9FN0SUg9MH1DlpzUZJZLKiACjC/Lu14YDz
wU3+Iq8FvqAfuYHpdT3tvKaeOux7KWehN0aokwAjlVEzlCIj0lEpRBwCTHoUS+O7
S7aeK6sv/uib2CYrC4xPS7YxjzX097+L+8q8XphYe36BDOIwf4YkgTkNn/gfYR+t
FuBziod70J82IlufcGm0AdcB2A2lIabcKaSfAh4bOcCz9/K297KArHNte/JU3KXf
YE5VfKVP5KN/jNRh6qz5LkOVhoyZ6XFjQ5JBH74G++hQtLRNZVNKYFtPGtbfm0FR
wxy+u57QkJzWpNXroD5WExxh6oT9zpEbHaP1dzvr/yd+7p9li2G/00xKbxczwNNH
CRPM7zwPjcu9HL200HiywuxznM/wl/4Fx16bFmcRfA0bUBi6zUYzXDowuiExQbtZ
L8Ip+abj/VDDQyA47+/9Ja1LONV3eD2pamLPMSvTzdGq9eIPJEw2ONWqLsFWY4Cj
Xw2g+HLxx7TUKznFtqoA4uIxULC4U9/V4yJ+18bvwTs2Rd29skpOSUf2Z2WO1saz
rZP+Mtb+fnP2yg8C6x0X/iTSgVXywtmsuqYQYTtoEfb3sDpgk8QxdWc01VyiwVah
NNLSjqW4KT+5uCxVzzWxMNn/pSdoD84X6oAhNb3bKBtA69p6wYMqEIIbsIaK2UyE
SHpf/gYiVqMLggWRfE8bDBODiMGSx9+i7JMCU/EiWa+JP40d/fPNnnJjYx2brq5/
uXEQ6sNRUgVxLg6k6NkRR448zzQwYyT2qDnz13MJqI9qDRe3C6UrBc512Bt4qZ0j
4pOyrGJjEjqr22zMfuSWXG9ecWJw26Liqb5YvfE+sNbCIafyDjc78dmsu9LmO7YD
9hMWX7TJebMSmuHZJdt+/jmzIwg7s3bbC+VP9RvAvE/6mTjDFb5t6yRG4IaQZX6H
buPxsVV26uCJCQYTCu0kWFE5PVTiBl7RNBjzCYcNlSMD9xOVOC/uOVAmIhk2ANgg
CgUOAk3CAwbhOw5pc95S6OtNBXkn2zyQ1qQkLNrogFR3dN87V8jHVhnVGgCYwURV
Q4yiS3ihZK5+xJ29JLJOmysAqerugFZxcWpGjMIQNSrtisPuQF8KRz/aG7G4a+sd
ML0TwHWbvvKRE8QuC6TgI1fxM0MjC+7f/PDxDMq5EJOqkwnMjyU+09WpmGkyyYCE
PJDhPJNPdfwPg6dHUbjBzuaZ54lvgC+2EvrTb9IqYlaz27irpZQOWTWOLRyzi9UU
gSDO2kB2hNw4T4iDxLmixaMwFnSXo5IgTDJ32x+VhgTgnpksOcA+gTRWWciQQx8m
Ee5xPgKk0aHcVSvWzM5lVWvobqbtZB+KqOso1wWaxccnQtbMJ6W+/JVVC7y8dKIx
7Erfvt/qDL/WxatQVPwNwM56nf64g1yGK/STQnHBP2ss1KgijqsGmLOR9aw/sUPi
METGRByFfn6V/iuJh74zwsfiqAOClIOyz3giWaDU+u6HvoYCCOV3lkHv4MXs8C2U
pkRAlUDIWvfs0Q0RoAX/GyR/yGFs2BoB9cJ9PqvCFUDKEpEhoOemptuDjANX9sKJ
k7SgcNQ++xQgAIhr7nYg9od8Mmagsk6rFD1q88ppYedcUnP3iXyG7Tiisk2XkuFz
J+m4y4k5u42MayubINFwrjnG0wAlw73v9v1bH5t27r0=
`protect END_PROTECTED
