`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NxT+kqYMFLxIpXiPbtSm+WLVnv3i0tpCjSjSc51YPLQwTY5VWLqb/AMFYsasHzrm
UquF09jintiekJshWtJlmYEp0CpoUYddTOF3/gKwSNvTnfp05DjaiA2n0PxrKuvG
r7cESJ5ghKN/QF2WhvjP4duEfS9+CPES9xlPP+FAJnWXxHo0InLSIlw4EgvFkBo2
064J8AYpyx/f6PpAEhO4+XwiSAQNtIbQXmXtMBjsUT1ux7Wbao/wmvYdl+KmkKiR
+NnXP5GglAngmeBmtGlnbw3AL7YRbBe+4MpposFevHbfuEFeZfg6JKnAzrdiBK67
LBNXf6jfNtRHQ5sk1o3gL/sHNQpduulkJJ2SxB9NT9DuM316tllotcd12VMKywEq
iVQ1zTmrlPeJR1es3l5znRlR7l5dVtJ1Kh3Ovvs4RFqcXwdqcGBKsEpDAGsrK7Ax
Ql7+/blE/12nIQSLVh6MD/R12Fn+DuJYKFkXZ5xgdEqczFaMtihHL6fmjzbnPOeF
Dc3TRpgxBAPKDpQ7I0r1JwIWsle6eOifY7ZWSTZQ5jqr1J9waMtBfzA20fJ6PwrF
hxxe9k/CXkcDK/eLDc8YBrWf6RHqZJfLhL31207vg2y93HF5Vw91dXE/IUnQkZaN
kxkg9TaUcm/QzfwqeUGPbZ73Sv0a6EfutYyATXQ5pBk72mlQDoF5h39Th6d6BCA2
mBs2ENAZXX+Kfn5askC5Q40huFgQtlL7wXN4EELFRZFH1pczDs1n8l840IJwN+T2
7DC+8iuhEJv8Bcn5O5ng/shBGuBVT7rZGh83Ol8iaXQ59Vvk/GhRmj3aTUTjqZew
Mrd12Tso996+pIz3jvg0qprahLn19McBafEzURfd91KfRujE3eDIOJwIN6dKByNq
EcVmqF3t/nujctq9nxux46Ku5WMVqD695RT33oNGaf3hzi4Q15PUyCuBvMO5Bc9N
tOzFQn89YK6Iv+tpsEizgq8G2o5iIgSl5iNcGyOXOiwBhlkGWRFW5ZfdYe+01NH2
KNU8mhAeneVf0XfrhreMsYa0jX8NaEUc17nnXHGBGo8BMIJJWO1OhH1CUImKAAFy
a7Kg7Fpg3AVJ83lObBk0SkS+xZogFCluRSvpKCRV3D1ypWXmz7eSLRcCHBAE2i9q
TS2USGrCcJS+upHvqBvQ5uPjg/HpV1tWN5E0UW4s90wigOGZ0+nu9+ntfQcVBW5G
XQI4fTEx8PORAUBsvQQ9ZrGboEP/+OQFP8AyEVX2rIuXxqDEO9YdnyBHwfsMzmfu
nYQKsUTMG/omja1omoug9NorUyZUoylixXIeyBN7knvlHX60OXqBJLtMcLJwbjYr
IgTrSlcIFRuIvbOC46vwS4m1n4i2mVU9Q3/Q4OdLXp9iLk6afDf8maDttCvAojZV
ShG0XtTOvEjdC1wEwnmQPKZgk/+I2fXjuPAx/HEJAzd2sIxTiSdX3y43P6d9kXzP
BU9+R0A++g9FYTPvzbbLYVlEx8x0H1d53Z0chLaows18IItyTRNxk2Frx3qvF++o
WfoaH9urY/b6zWF9eVPH4zEfUevbLi3Xc/sIWaEWo4M0Nl0Me5S0mrIVRY9Vq0X6
JtK7pGXEXDgKi7GqNZmNT7bU/sxBQmooNMZws15psLh8Gl+tD6jp4EwNggREZyfR
6PQEHPkJQuUAWN6ysuLQ9U45CVAMmYPyeA3PIg1kdHFVP8SVAGRq2oCmrjfp11mX
/zWj7/avXHfYWiQky6W3pso3bfiSn8znhJIy8dHLGvZVAYn2EFuDTmsP0hBVNsLV
OND9JHkqaZRxJWcgyTHu+8KN+uw5Pti6bMQYQseYjU/c2c1uOCvd/2f8exYGc4SN
pgMKnl2i4zUSNYD6sQJt2VXo8GQaAelglXOAqfo3ulrwI47Krxbl7OYtsyDzw9jR
+/3pDJZgKnOKZXkpKa4X51Vdzf9+CqwBcPHtLB4gj4RLJSYcMHUkCIvnlIpPGYnN
zAzvIAO1MPWAWpu9WyVlJqWmTa21jFmJ3T2dDH68dSoL7ceOpdYMYbn/UAWakcAZ
osOgOv7/z43Z69FUlGwT06/Wt01fO4Z1megXw8oHw/LmtlwJ2n3Wl8sXk0iUS4hx
czrfzDz8Zy1BdRMTPFh+gACtmVpWmjnejnuPmy5RNwrZPOb9LPIoOHynZLrvvUIx
9wHQZA+JovTkVdIU063Cykpaf9uw4SOaazKEPjWnade60XuOcJg1c97cj31PET4f
3GKFnQ7MD+HRPYSBBSbfPiiFVRA+EQDaBK5/yBMc/f+cxgAHZpaJRoSYbl8BaCXO
hDMrb1yAIQvcKZdEYusryv8Jxv3i33G6+sGrCVKFSN3KjWI2acRDPfT/ke8ckFB8
YwNrvT8LfTW25od5eKm5Fi+ZRtROvtdu4z9eKt2yGnwFmU/L4EplMqQR8BgGgWRv
FwOEPLkMGbw6vLMAc7bsMMzxWWT55nflivSAoERQdEt2uyVZsiNOuNffewRY/YYD
oAZcmG/NyQvApMOXmgvpZz43Q6OIVE4wvPCpwDEeca0O5GXzx7CyoJhZFCdjeYxC
EeScgGD3b2ATBkqqBbmXRfin4g6zYf0JBbRIgYkZGmhJPpeJJFuZrp2qaJjI5qJY
1LrMp3/wlkJlRGRmf5oxuqsFYKyBqooYpkt1PYMw29Yt5hk9HPDdz4NInCdDrSHX
IBunvCZigWPxUFY/H4DBeTK0f8Ia7WHzrDA9Hg2jKZDzWZYFCVf7LE9rlSS3nPRz
yPfNSNQI0/lglL4iOuHhpJKaugyBAiw5S5QBaksoV+p69MiWVeT8rpYpj3X9xf88
SNAKvle8RSwRd6Xy0rIw11nMNSYbdoHLWl3kUgs1W8lC3Z45s4YXI0zAmcoZLF7D
iY8a+h17deWy+03U+1rbHx/K5NhnP1U4FUoUldOihbVDE1C9Bg34XkIinnSexuiX
QtS05w1nkIHWEASEUX8fi37aSwr/I2TyUaikv3AiQxsXRbtLBRy/n5Zi0X52Nfyo
T5nFnQ9ajPlC7czDAa8HenoQ0QV38wEvcBqRVbacx2ohMINZr+FT9sqXnL9SPYfM
2R3qxgFc4531M+QuFIcl4k3dbm4sMVbPzfZEmger0eUofFYBe/vG/ETWWzlRCpGT
XLFHl7+Fs5gYQnraZjjZM9ZnpizvN4DKxWo0HhO48Ob/Qm3z02gXmnmzNrHr9hhi
0eHUJhF0qej3rMD6x8XtIqN2k7kf4zWtaE3wQc++/kRsjN/S5eOLEYqYBEuMoZsW
/8nswxzm0q3lDzESKghK5qc9xVdUVc5XSmnVDgW8atmJ6Gx/xDrJlRZtf+xG/tM+
72B1IWZOshsqjcglKUp5b8CJEzy3f+iDeuYmbnV+4j4RaOxeYRpK/DzJI/7SOesl
oTFYnAakKTiRJ+7QnHvDQsQkqhMMK+vNCRSNVWVR6GCgbK/kj1FqV9poB5YIHdeI
zIOWyn5ONNl40B1I+CsCcYYh404ae8XOoHXZBgHX8wdtKJtAC0+cOSus9oVMFGjD
HCKDIq83kaD5AqwEbQG6nc4QbuDSgWcrmLCUyvDtPyNXiEY1x6N/AtpvX87TOt5v
zoPb1FFFZJTboy/taR07t8PRhnVICliWFly6aQ2mdLghR0cSJOPjc9GAvExiJ3Z3
7xQomCmpfhB1vQ0w851Ikczg5DAEuUT2nyBWcdOQlpOeM8+DN2q8infzlmuLQK3D
qYfHFfX36Gh47DhtuVYwURCwca+PjULmIxmbYc1jUu+YbVuF98HkO0GsDSx6c9i6
GeD2/w5ugcsWdYGdih3cc54d5b4VfADTI8raola5R6+YTGyLizMng6vvKmmk68Y4
WD5AGB97n58BQOK/5KSl7HU1Ok1lvopoTAH7/SC/E97GxQ2NYiXulnnX9E/J6r09
49boelVJZZXfpxVI9ETVn5MgHDFs8fVWxEHHY045CnKnnY9wawX9u85jwXmhbAjQ
aQlJN/gRDdHr35vvvBZiJIx7NOMTtzJAt1iqQubvRnjWnU7ob/pUtMcpoYc/WwJP
D9J+VMETPiegBc/+VixV99u6vPvExviTCwO/71KOB7i9H0nyk6hMRK9e7jawx78Z
R3OyOunDgcgDuYL8JkOewQKTheMLxMT87RQCXYftLRZ0QTMsJhVjk9megPLku2c/
8DHbxOmx3cZuci9CXkQnyC3MqzY1+MiIEIcvFJ4Xk6rYiKPJTGBLmI6oxbkUGEve
e8ug5ja9rGCtVkkosD6Vmz++BDvdQz+1nivaynirQFZj9BZqC10PD5tP2HDjxbEq
wGZBUYNlVimOrSpy5NEkRdoU3C23uwhnyWuzrwrV4jEc58rYHD87eMnQBoybZABf
cdEc/uyB8Zuoew44T280vloHBRqPNvsoo8fkcHVd6Xe8VdOL62nqMTdjMFbtl9CI
XHLQHgcKD3V0BLBl3YWyu9hnzrowzWIkhdXiqsipgyvwDS8jkZbdieyR4dnQnWfo
L7jQ4YhCW1ACEr4pgwSmhwEFju4tCBZCXQF0hb+2hKctKZJzMAJ15ySaHMvmQIu4
oSKYRCIO3/8vvIafdPp9isTAOWz1Bi5a3CnoV9uVis2mGcu1YA7m1w6prM4Q8Ea6
aEn9WlR2lDNQxj/5JzyQdH8GAac2b+FCCZCWdqUwguo8PPDwcxFw9XVHps3Fpg9X
4ISsnRXBaBPH3ySepHCCOMAFRG0mHwuF0xMy5eELVi1ZCdomWQYvTD6wJUJmSbwC
TFxsfbXqzWl9aGzDwvJ31oyjZPQ1h4BH2jftz3vXNKio2pCa8lK0dOFHBAf1JcS8
Cn0NclA0z0jshXIhBBdWDM2ahV1eJ7qgPhPhtojnBYPrPogq4yE0CprWAT5VMjh0
CgafKa88sp1TXgDS9eEqMrUJZ7QhT2nIjTeJohNiSP8mTjBA3a9OkKnAjykt+TW8
Uaymt1/Yx5RRkV4Cmq6u+g4X8y6MispzdzNJvL0DyxkdxdyjtvCDAeGBFKyxgvix
YS82ATECCGUxyDaAIddpVK9mcIDW9Ykcf66MJS9x8fABGZKk9XxMP5Te20ajWamt
WIRTolYNfN454cYdjBkug1v6xA1K7pD2WUefNvTL3PQvAKf5n5NdNgMeqaMWOk/I
PLpE+6sCkRnOHxw6UKpkbfNv0m0yG1/xFdz06xtjZYopslMltN9SVz4jnd8rs8Zp
Rn/yRh6CNAVvx+m0yI6ySgQ1SO2e/SJHhT251uW04REXOvQYJO+yg5cVtq5cm3pN
HfWUwuVUB17AudliAYykcz0ywBvv24e/xzXJX73qafRM7DQAewRpxKqJhjyINwx/
Tth3sPJl8VUJJmpOPl2ijA+rjDoDhwekz3Y45ZST1c+ia8k1DLYI1lF9XhqKw7Gx
S0jmDQ0U4WzxbkROAKf565+PuFBJ7EPunFHvMuPz5qtT4RAlc2Ire3WPEkL0t+Kt
415SlhmDeOQsxj6TlR6XdY5RBVgbuaU1SWIq5+3gbNCMr1nyZiiRyFA7Wc1NZA2V
5tHa+BOCTV6VZjLP+FETz7TVPob+wmo2Of/TaUAMviTZy4TtZ1mEAVxTRd+SLCLi
sxcSfDVBHgjgwNKEPQwIRXDBizidnG1NKdJn55etT3cK0s9EQWbPOlNktRaMff4l
8X5Wd69iiusyBYmwmeCLZvm0u9RrBEIsKQ5asS6/KNi9BaobpJUMVEemYFRYaAsM
`protect END_PROTECTED
