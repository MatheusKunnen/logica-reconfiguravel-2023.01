`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DSPuFAPdasEK6lO6DRsq++P8gQkqbYIuMSVBDpXq0MrGUefgydQiIFmiOeWSRtmf
ELsL3H1qWRcCY3LjLLVns8U6IoxE4F4BwTE5J3/ReO7iwV2GTnEBK4S9m/lN73R1
oYpRjB4KjznDOmASe47vlB9Bt836ZtNxS7Ls7MuJbS9BzzydoEvaz11IsgjotDfx
ZDaKjjOkqZKB34Sj2J/mBFM/wAvIYueuD6ZCkfSQNWzYdKAziwii4eYEP1a8OaaK
6msjyBrBC5z4dcglCdRxKF2MQlIeTlgU4tlAmvLvcjdy+/451jzIYxEOsk8BOLEF
NLe5k8dCGVHP39WYDpAVhRgAK2oaUH5c+3BOrxmzXKSXKCsDrLwx7/3ClCGvgesE
9GdUkYZrnJT7Qm9U1cqq3cpjdqnlLp/TnsrxgsLZY1MoLxb3PJJk+ZTVLn215KG5
xP7Pwruj0l2Gbntf/vaDyeNCvh9qRoidZ3xqpTAuJf/Q8z/So50FH7XkVYFJbUyx
JOgVNbG1vjSW8Rdul61FRjJYmKA/OV2SXDb3nEoOMVlmqj174a3fTz73Rx//1IXW
7kGyzf2Zzk83VmobNwPNXal1giAWpR8Sejq03vEOrToRAUb+0waeKhYGR+Ybq4zV
HKNAdsbCsQ+J7xRGxevRhhTqwfsPL7L8Fn0EAsjIyaUPKMNsGKbRpTc32aIYDJry
z/hWXSLUgiSF0ibN4yH2JqBY1apTBW2bm0IuRs3xGilhHEP6Mw8y7UHavYacflwP
3ZA+lPwnLe0CIC3FC1etJeozhWC9mSxdUIw9HjQ+qm2KL+vQI6McqjcYdEObtd/F
6mOKMYOexI3DPhjXMkECCqJKNiA4XdNeVJJSYMRrD3qz64GK4X5keUCL6Fvk4a2V
21yTgaANN7bAEn7kvYuhd5/bqYm9weUaNes4moDkA6o7KBhXxCS+rLQJJA4k8FQi
9B9MRLi2laMjpaYKAb2gYaG8EXw/PoNiI45hY2bEVhNqQEy28oRJYvMrlxz9Fi4S
QBQk3b6cyzK8UocBEEPf07U+U/2kADr9GaLvtdImq+9O+Sc9LUgbpVG55Kc+E2Jn
kzQBfWA6mDd1I9ttMBzAQdjds/GS6vjKM0mhxxmdO4tCcrWQ3onfsikDRjZUoZD9
nZpGqduv+SvDxnkrn4uP6Q0H8JHqbJqjuGHRvtSdBJXkXlgTNF5sRF9IEWdAR9tx
o3MacLCF+bL6vbbfGkVT1uEruIOwncDMDW47xp7t9qqJGQC5aO1Y7lKCJDnbShNq
sw2i4rPCQDgWlEtH7jPW4gSZtU4ptlEedyEH6pUHPQJeV6FWhOBajUyNHKW6X7+E
+D3q0GSs6CppGWqMbEijVcXbP3oqfnZHyqApLTD4doj3OaP/LZCQkPIxpgOIIJX9
0Fdv6QI142jQP+LQmiRuJtq5KSJlC26KubFKkF4Pa3APtVg+dqJj6Vncn0mNYd2L
ltaPLc8xDLFUB9RAq4fQHjPzRYjQ19uU145ZgBAv7zCKFthx3S4CHzJ9i33KvbMR
nB3Hjj6SCEAGpQOArvktXapgCVMHqoHG1aVsxO7KeSnKVYg5ccenuQrN0hCRGyQC
4CGEKNZQtmPz6WcjqXVpI7M9iWkq2bMkQZQVMclSjSRLbDcCl8GBzmbeTe0/Zg7g
NnDOixmpYg0Wt+B7A4VNWsu2RE99FOn/Oufp3G4shKSI2f+mLiXRW8xJEAcptxeE
SE1M/3otB0JStOcbiaaTWURmuwjnHD6sMUqQPWABzjOfJF0Rx38ZnNJIqS6YhSll
Aupb56OVE0u/cz8z3HHbUY3/LCY1MKDlPQjZiCJTkyb8rj1x54XOR7Z0MBGUU02C
xiUvXgrlOB4qwM5J8iAKsmsCWA7oGwkmDN/UM1KqSMBYOvuZ9Ul6tjm8y4wZitMG
DoeTto18s1HZRyhHYieavHm8jE/SF2Aow3/RNyAq75V4lHbb1XGnMk6zf3vLCQjr
dotpSFp1YbGt/Ep34jgen7sdntXbxsSeTK3AhgzNTAGD5Kvtb59AShHcytpLuk/U
`protect END_PROTECTED
