`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bTRrKY0wck6Ei40CnVk8JqOucW8X+ktmPSBAY1QuVGCOOgb31xAu06ptX9v1OGsH
v2v+qkc5xGF1oBNJVmhsVZAP7njzPAwYFgZYZfhzJJZJwt882PpYqg8uetl7k+Y1
suMyNaO5dudwQyqS6qK/hWSfFgwIByEW9VyS2xMHbYH2DuyrT0F/troBkO30zM7m
0h7hAA+U3jzzquaMTQRCtFHERuMu40XLQnaPd6L+gO1TCNd/MMs/+kYTB9TTWKGH
a+LMr1FwoTCFV0W27xav8V5v1h231tHPFvm4akGsZNzBcYVyU4W3h24Nc0bLpLCI
ZqPN5aMoWLG20JPkBMZ0cGp6tk7BJbiWiiKAMUlu/EknfhIBdTPoLXzk9Q5iCLDU
eJ0YLDWw24gNIRytrCFwcJplzXPGiEt+d7kTJDfTXL1acHK84pAgupVjD4sL+cSS
0kTrHUvDYrau9ML3h7XJ9d9Jv2nL591IYxRZPkTVCCg1iqZvX6kONLtf+b+tqrtL
f/KavHlZhPRm0kfW6aEyiQ7fWaksbwGkB0Rcym6Nnfs6z6883pwrbN+60fAq4xfd
XfC2i/Drnu8WSEpa4UqXod4+cuQCDHcteo1mBzdoBgU=
`protect END_PROTECTED
