`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SkVVid2iXFnsCCS/XfJ9qadVmH7uBGvhvuRNTEX4W0tGfwvNk+jObAErhO00iZvA
BPDFZCrMuanPpFFXVNJMojoZZQxapAd+ybYhY8JCDQCUeSmKtpE4OVTn3//0WHgb
0HHjWTDIDvwxQMPMMi6ao2JZfxPwf9IrKTP7Rh8/F3pc1u7i+vz91rwcVBTIgmsx
ihm6EId3LqUHgT9/Q+KdW3dlH0hq2auF3xEDctnjunXYH6Zg3EtBDeq2Xd9kXvUc
JVt9TIuTrQfx1NGloXWWeB6iUafjm7xONpvgUyWCCn5Jc+GDFygoynNhrb89jDaJ
U42ESICPHSNIRSKE8wOAxudjxpPtUc4ijOkr/wsWBKamtFkmFGV5aYf1xhgCwBV/
1NpqxgvnNtq/5VHCETwwa5MmPpbYvD47Op5kCVije4XTcJUg7EFfshqK69379OQV
KC1VY5e6REe7LregnI9PFmPKBSy3/KUdWOrSCvloaoWs+SfCNOf3A9Fln1/LeL0y
aGuyZfH6MRfwECBiVScjBCubUpDq6qA47xNQaPn2s2NuYNsGWFerMr0afwQmiAUv
PkpmmTih7cV5+RIKE8HoJwlBot4/kXOfEhM+TXMsLdu9Sw3SaAtsq/sC71NDzZ8o
WeiFi+izRGQAyStAahNIkCFsUVGb7hwYgqgUnK1w7Z5uPopxHoa6BMhx/8DMEZtn
jhpGXxIabTUa9EZAtDkO8mJ0fdqhkRiZHd7t/TET9ZSSYE4uvrL6Xm6S/bd1dYzL
KUXG45i0AOzgAyTa5UaRUWVm1h0uJppfOZ3FhS/c87t1a6vRqku3yL2ER4leKu+u
7rFYl9A3dJq1kXJfcCCfknU3MUXO0BRr9wwF5r4giZQ/GFCDUm1j58zz9cE4A/23
V/hiOFlWdprTiKLf73Kq8KlPMZTWFRMy7Mch13Mq+dE8Kw2qnhLo6wVCn79hcvBb
zDGEBKZWKgCMQCMAPjDkKCQwsH++nNvmwZUJjIf+OMOpocK/200+bDIiVNdmgb9M
JvmseMOmWVocvAEWIOs12UqUninbd7FS1qHYr9eLKWr+tRCQEqEJ6W3SfQ+BU0Tx
ssP7cVg2+eXJQJ3fpa0GrrQgsPIgp7kHz75PZ6LzVLCl+80uvG36ud1KDb/BM6Sh
6NO77rjJE85LRTDHClEdqULzfth3GE7qVpO/B9NOdTSmGnjP8cAE1e+HlYMn+HRJ
j6E7PqwvbvWdRSfFjghghEw5QaCh+8z02+Odxkp24KoAPE0GXKaQB0Lk5LVKdi7I
4yWHO9l8X07aAhYgewtfk5NyfvsYyZebi5rFkaNfJe+r+OSnl3X6bUutuVajq/Qa
CLbGDaiUZfDrnp7UvEGqmwPfwzaQxaboIr3JrGk5QvKkGQmA+derNZTEs8aIDdD2
ERinVeF9gfm0CtjByS51WUe7XgecrAGqXY8hpYozDvMBJh1QWuOcM7dS7B1PTwpf
y912QkocPNWJdAM8XvpBXHDkpr2do6FAzpACqsROFo4aIU+q1hKIvBzurIJmBFIh
ihuHoUMiyHYDm05qB0rua3atOGP47gd5kFrufTeAyG4/t938x8XlkZUUg+M/8FKJ
m5t6vrGRjKrhjcE164v3KTHTTm20WB0EEUjGlPGrhpiopgx498BjDNcRSLkpVG7e
nR3wE2vKLBudMt88aF2nQbZCNgoPFiyih0Nj7FwSJ9BOaWoVpqmajPyD1EF7M+v+
SastNZorZztMCGAKMf8N+Irc0RfhVB5Ih7oST3JvyWVv7X3kLK0Fmn8jSNjc35Wa
HJJq4gHrGtlWGDwUfe+7rhP5W1Kc/PkEGMAFffom3vx7meXHnmNiJdTzyYGWnhx/
t8/NkDb3CopQ5Xd3Uy1sQtiD8oajqJ/C+yai1eHzjWfrbUn2g9iMAnGJwtA9B5rq
/0fh885Ev8HEHovHGVcoeAQWoeICh94cuY34KtarcOry9u0rIKvMcpHkoYo/dEma
VmneiRouIgdtz5alFl2iwP0vUSmilt7NuXPaGNy/arN9k8TgAkVVMebDMD5f0wrw
tTtXZ2bAFoC/X0amDToGMg==
`protect END_PROTECTED
