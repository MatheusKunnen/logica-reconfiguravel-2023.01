`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VdlBslFi8F5Ce2TwkHNq9qQFnMRt1BPXxRwbuTSaSnDDBTTzqRefWXMF9g2jON2C
CZrmeR3LvntVqj8fs0C2OaJcu0jJwFcEbUvry4fFHSBBFOLepM4Gpahl4Va4x2O7
Bieu9gM9/a62vqM9QVRLWu3A4m1Ys3WelT8NzVcbPTcZRh5cPP/pABuI7/0PrLr8
lv2Ni/76iLWGWy67qIpBJwcSfOvhmxgcAdZJMTtUyqsQtrOvM+Vj5IpmNljIuvFX
TOh+CrE1MbqXGVshEzI+w+EUsgBQ6OYztznvbm09190L4aZ6JgwX5uWwAsbrK7kR
v/fYG1fq8B9iOdLJkCM+SryVuwq4NgVTjDsSzmhsZajST84FmdYswA+xgMWsBWlN
2imT+XImkVkbgDTcf4EEIi5AYGxMWtQy3yHJpO3dlBVjFpBpzEGO+bjQlel/FoV0
JXuJT7yI2tPHMB5p/hhmejQWv8S1TyzneCuptoH9ArPYKr3CO1ZQR0mUpCKoobKp
jcmBwq6wchEFDI9eNeHdei5rWLTv1XkAe8/xA9ur8hhWiAzdYWBjcmdFXT+EtLbg
3P9vLFZBQdF9IpuYC9Tb1MfUyQuNpPWt+eclZrrw19H3KNOXWV0mrZz7SWR18Det
j2GYyzlImy603HqnN1fnrDzV9eWbSHPplblt5Q2dUraIzN6k/Emh0Zk+cQ8N+kUz
hbzYuoG7clK3rbtSyf0I2MwIfZxapSRTVmyi4HVtzb5DZhT2cAHN7G6W6LGXLL83
HvDyb1pBlbha3+ZAJ2RssJxs4nIrQdOtnYpgQ5fO2cJ3OJRgmyDj7NIFNahWQIlX
9I+5suRgRFQnlEhelcWXcMUDOjw79cuHoG7GTyzJUk4AkV9AuP0fv3Pt79bNPuLo
EwpUVwIUYJe/eJR8evsbIpFSKXdJiUp9XUWaqzgMRpWvpCHE5AWT2T1e4gK0eetX
6GXcfr/DWqpL8VONmjotwkEE5S/qZ8/gyNUEj0/UIHMPL4t24UDoPkHTimXk4DcH
3NhVVZ2jqwsE2OVAQLGTdBgcxNlXeWEI3HwPRH7q4XrqjdnSRLJqLsFufwI4hd7V
OwJOUEh3z8V53oHaVOKPVnOG4VXSTjWbyfSVlaf74FYGgy1mkhSKAT2FHMU01Qpo
0cLyEATbA4ADK5UqMqJrxSOA8RILcu2uC2qaa4vjE2d4UbhvTt97tOhzVUn6qZXs
CrzYSpD3dkXXytwSGrmsdT+peH8Qiig7etsaUNcbUqP562QsSjzpf87mDZ6Tq1yQ
u1HwUiUDva+IICSl+qPSjsCakbQHdcDyqBx8EKTYerJN+laTQoHL//0/L+1/bTcd
oB/LqPURgBsMVvlEhtUtwFJdAU4tI72E5eDVe/n1weLIdVgyl9n3zuK0tddeY9ou
NTNDKp5FvOfNSlLrv1y4XscQDfkelHK8A2h/sDIB2ZY8smMOwZCTL0EFI9eQQn+N
FjJ6/P14w5lvf8Ofb7xQqYcB6xoKFzNcpfDlJhLpTP1+c+I5GYENfLIILJyi2s2Z
/LhuFWBGpCnJqXD4u5o6k9etrqeOyPr8MUXoWB2HUqfFf4pnFoq/N69Dv6ZlB74i
r1ReHDAudMU5YBqX7FRsmr1VLcTbZkpqnEKkYh31op425Yu3YkrByoCd6ir3C8pn
RMtb5TLmMZPf6n3m4/iAWPQKAEau5YzTL8p7rFpgTZbOkY0plyQFqeXZzaDzeLMo
gSLGAFoWBW/DB/86DrRbBkwJjgRXYeJ4OS1Wxk58QvqNAeoGLWEUgS8fueVNH+Zm
HaYZn9mVf0NnhWrqu9xLN2gZs/7VDdyvP+VEXKKpDtAOkm4P5e1YR+dw0oboKxcD
va7QHQn2c9Ksb83KcniNLNytR4f/P+Sb0LiqhcZIeZjJKnQqA6gNtCsov30r74Nv
96Gf5K8/Jo7tEdubvt6bO8tb+oguJqIK0RhwMKIaKufrZqKjHSR98km/aY4fVpj4
RDdZh7yDGFKZ7MlLOo2yhYrFDv/TPTOokQKrsFM4gWcqGe+GeYGU4V9bsDUlQq7i
ZZR/bHq/odnit5GLoXnKElKQuzBsB8prTOOylVJ9z0q+JXhXzuYwr41IF/VLow18
B+E5pJHcw5dSD4w6pKsZ6BG0shTpPnXNL+uFlScLWYByI36//mf8tCR4R+xAvo9q
6EAV/8+1ec/ZbFlo9BA4yZlYtx63BlYtjMlko1BFlSoA8vHX2V0MplQM7gxRYroe
d+k6glfTx0F0kxAXjCIffoBky+rAFfZIjf7q5pl0mIyimFE5Pw5zAa1iCUgNM6Ti
5/wT6A8DvJ9grukgF1Fsy1nFHMs+uatZbSh+NZiNrD5yBA694VDy8kHnaCHhEx4f
FxpVMPzmFc9UFBspYshGzvLU9i8u60EhtgZDRnas9TiafmhwEo39B2Zzkv4v1Nzv
FdYsWtahhn5vG/rZK7XZyCYOqaZ2iBp3pr8ZTYTgjEgyh38po0JRbvwWb+33QcKF
Q4FknxzuX84/BLtDO/20NMPTKoDtTJyI9WwK1USFrywTH66aEdGky9QOqlGhF5EU
g9/siygezlEdaS51ydBslCeSB4ue01tpbqxWjVxU97bD5Sz592W7avNFNdDwguZn
g+qnrUeE8kXK0ggQ/zGlqnm7pSUIVbe+xHy2u98rTjUPUQz/HLeGjEoQlszbAqjp
xgk6I4H9KwV2QmB7lEq8vYjX90m5BLEEOrNJN0TqTEEu/HUyBu11I5YqgSm9WbY0
/y1zsFie2dUw7pL2GX998oxinYnX46EMKD9nX/PI0t2ZykDwSWE5gtw0gaa/Dh0S
qNm/MtECMGWdVmsXRoo5Tep5GREa15FqKwzBbr13l27ZgVqjoXB9Lzg8t9oidcva
0IPRcraSfwc4VdwjrMsXA8mOoVc5nMfW6gONY2xYNIkQZh1BwYnYh+jX/45/181g
+9aN/BhFHUzHjARAUP2H5+G3k7vKIq24A1R2Ga9GxzQoFoiP0SP1qJMwULE2wCDG
/8zqTfJ7NfiXtCvCoROlv/EpU8t+1NoFf8lnsj/ncaVSK6F/fn1sPhusfUiSeIAI
szECwDwy6dBoScEOvy4dWYu6yfYPHsTsSA0O5zWBqgvZjzhg6Rrxv2O3tAnnUHMZ
4qbMsH4VP5QvyariJNeDl9+frv+shUUo5CKZDGL2Eb29Spqw2z/6/xsTukv01l7n
Y3dvN6fVW1h5c3HSlKd2ZBz+AH3oSRlhxEAfMGlZZ5WhPkFQj7CPCDQ0JfXMLZCW
nYgh4h1vMNizhdzJnkLXOc09L6q8hsKKYsa8mrotgs/RmdYof9V32McWvzs4GCNJ
J2xvMKmfIXf8Irz6Tf82MJRSAUVfAdmQPZZmBzThNdKMhA1KsjjeyiRH5HC4MyOY
/5QcyJzXM9IVrZlTrMCd26fQhXojQZS+5ZrCNHdCL88OCHQc9+ZxYTBZ5PwUNCbH
DQiLGMpPOtkSL5UaZHtOvUKkEyGhyUBGVKwcUOgqs6kDdP9j0HQXmoIUangZPLxE
DC5XFTVy/RfCcwScklHhB6Vi5cYubJ8mV1/6hoX2TTv1+kubw563XJ2TqJ/g2JVM
FXRHFEEbl6Ct4UJv/TJzxLwdb+xQD1jYURcHSbHtalBy0YmGbPdwAREQP84FpFq0
G/Ld/J5Hq11Nc+ym/1gxSCOZt58y0mVBahx2KiPzdA7F/vSEmrFTd66PY9bJUp5k
RcUchjUYVCzRHuMQseUc7XfTaSlBWxmllsfeqj+UwuoQp79aUMajMgsNUZfR3GH9
1303V89WrilqgodpvywkQ0sWxsqV0zDMmbasCWaQnLQbPGSTP1+vH+u2t8UUDESo
qUtc9DaE6YmFkfS7hprv3ztm9ULdUD696VNdd5CeFA3l4/8hpbVsEYrmPJNURLDf
AkSVQpYHrWEEenDEsAt23b+H4vgRqTgf8KfyEgdcnmnpm13ZidXRbHt28dMMLNzi
cyF904VfYx8Wt9R75l4ErWWzhmJYtBhsRAQdU/Nd9sOWEOeIf4o8ILekDN+9DEq1
c8fgRAjT6C8g5B7XhBC/KZdMdntChpHmF143LPGScmDKUCAynqS86LS867aaQWpi
zGPGJAB6T1VCRZ3qRwQU6jMSaUi8qHAOWVrx5ZWKVIu31keTV82C3H2+GrF8ypxi
jRy9ApEql8AITk1CSeYh60tsv0Zg1i3/YKeiQj0cfEpB3UXTCbdN+WfALO6TysSG
Jdu7muIgozPn4Q2xBs0BFCNJj++L8OLClD5U8fT1Ecc53H/ESB4bBysQP/UqQvgv
/j/49pT0x27kyNINnzoaTlk3GlMwPc1ShU+Lvzr/OhEa+StaYf6TcbGUB7iG+R4h
2zdoJHNxztk/5KbQU7hjOe+tTHTKDPzB0HM7RCjOdcEm8SXDcV6BNS2R6TGBFLEq
cRmJI/h9o2mHpRh6RJvJi7tSffIlWwwMNrY5EtVE9eAOZ8D76If5xZ8yAfXoN4yG
hgxNMNU74yUjVgWZ0G3d7Pqy683+Zk2Z1un4USeAd0aAq1DOq/BaaIlECIpLIFPV
MTCbYmjmLIliEZW1YS08Kla0uDZS/BR6mBdCvccZoexr6hTgykeItPMZ/0YzwrMw
lALDYoN6De8Le9/j7fEaMRPf6By/e/UXW3+NsPmam2SHT6b3hMiESzFTzlSCMRQw
Ng/vNCf7ksLpv2ILr/vpUXKMLqMJ/CbIZbFHqClUUgosaXoI59IYku7MA9Y/I2sF
pCK68kEolS4+87WyacZPBw6d8sj4MMMHTlRtA3Um8A4ynTI0gggZr1v7MBJI8O8O
u28/tgfeGLjTUn6FBtYh9VQoODLYBqesBGemHHIITDEc2j156a0OdkbdnnSUK79y
4FomBuM/4BC3fLF45dgR2JEtTVOMmqIXjOY2ihwgem9wxDEoEZwy8rSFTguVR+U7
rO+9lZNm8slkmWDdAWkAQ5abKowQeLT787k4UPRNDyGbixuDJEiMungL8ZrJucAJ
h3jCYBYu5mRm9WsilbXN5JmkSz3cJQkFOLy8/nA7ML2KgzG+gLDSk1mhGgz+WrqQ
gQxCwwfD/Hqn7INH1cReBdXaUUhrhe6wRKIVIIqzBq4JAXg+J/UvnuBsviLqY/FR
Bsw76xKb5ujW5UjEdOrPsQX/mrgNTY7rcvGy/I3oygEQhpJpKQnYHRkcrNUN/EWW
S7pNLl784pGlgShXSZaoTVwQt4fdcJWC+RmBJX3l5X1+bDknv10+1cYwlXSEX/yd
rx5AcAm12UOGth35M7JzVTvRJWauWojK6eKUfOVg4++fkBOGzO4RQ0/vrk34WHWp
PxV/WOctSWXvtMQMiXlzdaV3295R4Qvkvw2RhhLkCpBU4+GCuoobUkprPTTDoMx2
qHuS18ygpiSlqLsBoRZ//CXxv0a9Vf97/IfHafu7vNcgwsecpLdcbUzPrvx7HUn3
uZoHKb1cxEjTtMIbUPUTnIO0EEzt4QqrMMU1bCCC/aWBk2/T88KNVMVFGdSOky8c
KSca8NZ3dyU21zgcC+MOx6SoBCohZZEgM1foBuoDjUVT5EoYPW+rEvkCHbqMNVny
LN3cA8ZD5u4s9JvmPdq8FYadc/Knh0EuJyX/qjTWWE7JBzs94gv+cfo6PVub9JqS
U1cTAZWnyJIuE29+NYDh4cVj+upu1Eqh/OGGXd1mqV2xYxqDbQI3we17QJ9aqbpQ
iKVCZwfu+kPtrTdwonXRv9MIvBZuFvsIvt7yVPAcCTsVuK4pkviVJRlGkoIEmr4f
EsxCAj+z4kB2Qd2qg7uTwhAd7TYzgMTQQJIwfjye6VPNJzfoEui6vdzPhyuhVs4c
xDsvilT+DFDzterYuQfot12/BWqyAyUrzujrrh/j0Uks2pQFb0w/aQaHF6BcE8xZ
ub6d36uYZmjXsXa2+iBNlQFFKI3CeUbzYmENK/0tufk4r3f144XkKq8x/RnlpFMw
9+p1KVnwrL1clVatrlnF8R0Oolf7LhKkPYdXONfUgJoCD0ByFolXqarcvUnhzBAx
4H6Q7dt7al9Jurnw8S9dVy1qIyrNAJFiWUvF7IvTLwu3hOowP11uFc8bnEda8mMw
oNu2Ho8GMHvm/mcpa52xFxlV+PeLEWhREMPPNkf54vn3541idrGRCoanG0nU/ilp
b/pGzhU4qiu0qRckVSbx+4Loqq+8lVFJIHtmFffapoF7zgVwAaUVwKy08lzH/gdr
Q7Eh2oAECe9b6VTqKPY9nciI+9ITEcKl/IfmCP3lqMbLbCsU0EZidUiYkrlGKzwS
1HJLwY0NS5D1t7w41tQoRt4tzifteBvofTSmDUmbPe60cN6/z3NBvHXnFU2oK03U
TDguKTu338+cJ1mi6zLHEcVOk61Fl7AXmvFYjSph7i5RdAMBMAR9GONaaxHviIUn
mwOuDycY2DjkmgbKwHcC+4yL9JHxharLVl6mnxH3PrywP67sXRNhpZtrbOrqtEVs
V5rfhd5puGufONrxHGhrzgs/RDccKO0Ygr6SjvsW5UULXhOFoUeQYq4387a5BviW
9Fb8/TOIIQEu8IUvTslJd/wXyZGOGu9dx3Ix1LKtd6CTg/I4V2ludhrvpJTMImwn
fH7IY0foaaTQCBAzGcKSCusBLYOhzc4ahyCq22Ow1sjfl51Lkktz33xK9z79AgaL
nY4VYDhW8vlgjHMXlH508EC/GdYZBLOeIaLrXgS9H91MCJOFvy7cewFYf4jqjVCn
bvqbo76ENh9+w5EBoHNoP1AK2MQKvX6c8yC5ARCwZgJ4Qd4iUl539Xl/HiQjLxDz
7Mik3r+sLR7bGFAzx8XIUFaaD9lXlxEWGcpoPsLcd+Ksfe6UEZIgHDCvboQxwoK5
yfc1w/9jjhPsSRdlsr7r4/C4CyLmdbn+9171Jy4NACYIFLgj3UYBS9ghbYsY63IY
1YW6SzXQZSm3WfsKwiiwFz0V4L59ymHUlIHX27RE+Mv7UrpoShzGBotPEStkk6vk
0dSHoDyxDTaOvHXhwup53eAe1ZF+i6upQEz5fXgc0140VLrC+eY7ZrmeLPuyX+GB
RfcqkScxn4R0PlVhOCOWX+s/YPCGGU0J5Mj2q25GnYIoU2sYAzoZmsnrhS0OlZMf
6SdC3opAQxNk+fc55Jd1FmDxO7zAxKG/28MQ0/+k4RSq7sl2VgFA5CE8FIJST4EB
KtJTEfguZ5D0XVHwNL/avqxsRfhACDthEMh+wT8ENXLa0NXTVY+YY3zB7vqV5sIL
2e4CKorR5ioE5pMIWU8kCR8qEbAJaNeVuj08+pjuJYfsJhQLetw1NDtwqZhRLqir
GT1VRnFjn9R+dVnXaYY7ppLbfGVQuP/mB3Q5y7M1fXD/Z7954tXNICxFg4HrYxRj
T569uh5q/rnEpdc6L0DRCEgDX4CtcmfyEmpSoF3bBvskxza5NDV8nNqESMpIXQLx
hXz4UwvsQKginvg92hWah39wkyoH7UVQc/M4Ff9FebLroaDbgqSbWEtYwTWKcewo
RyptVLsR91LkadurCxh9gOtJIiGZXND0OU/2Got9zHWMj4Ljdgdk66t8UIMDVTow
RpGqC21Q54Gko0zGdqTrQ4VbUS1Whe+aPLwVo1eVdO5iNXN5qiNec0o9oRP18AN1
ZYT25PN+1Ue+jp9+D3CBINaLV0URbiukZmt8NsdkOEpJDYana7jzcVEOaj+/gXwQ
`protect END_PROTECTED
