`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EzBTRxL3SSFEtPO4c1brcJm4JsoIBcHNLeFdc3hfhPy/5A6gADsAdPOvF4XipDGK
UjPa1xA/6JOIIsK2muKNzMBPcQcxaPl3BLOjOUU2I4FFdPhmhggpN0zc7htiVB6U
p6FibkHTKCGU66Sy/Z/h/qoe/1TPthV7f/NajBA77qUaubHu63cMsZVNFRpq3QeV
g1PrNkse/ersQmEXSNNhZ+ALIIc5CJO87gbuj2N/ignuRbVIKkE4u8C6LJ0I68Hm
vCabMBPCzYLvDmqWfdLwTTIi6Jxz7R5FEkX3RCNsw70bvtW4cpeGGt3JfmtCvTan
UMaqcbIC0ewv6on74QaRwbDkhDT85Au7Hj2ISeUVxnrdEs8hl3D0rOOj2r2xHDV7
deBSLX4m/XxtePqlpXtBluSWqfW4huN1wIrmzNFZcUkK22mGWqVpErd8Lb8n1asr
gbRI3l/6LwWbNWIHOX9V7Hw/w0YLcnkEMlig/JiVI9cC0A9W5+I36OXpNn0Wi2v/
lsoPVjUfdtaehTjcFMFTBK6DpaInfMn8q8ID0I12BRT3ACmGDS1GAtFvFhER8Ghh
3hFj4GtuX9ixaisSSYpQwW9Tlg/FxN7T73JoQ8jxB9Q1GbkdnsCQ3iY2mhlTFqJX
Uopzp93gzQR9Us51u/4mLCx5d/wBFc91kFhasyVRxyCxTxFIloJe8tzady4cB+Ru
REE6kLARohL6Ov1acr6pEix9YKuQftsts/s9nQ4DGXvAd9LlkgfPOOgw5A6h8XNo
mn5lIDk6u+vFuwo1wYFt+r5ga/7XnIc64i4dYuW+AF17lG1ZS1CQQYJxf8qpY3Ua
mkjM/QjIhSuTxyk7ubl7JUehR5Zjn3Pud7ZGEWKMxghClr1MrJ8EBgp2kU3o3v+X
stzR0bx/dwyQsIz3wLsLpjcfKG5JLAbLR6F/gDIu6QI9OOAG5YVcGKzudtuTRjFO
7Xqn9l7hGBJAceovwTnjJVBZU94vDX9rsgWyKJJfdXYJXepVmZjXBOmSyP+ezf6l
3VDBZXZ/4tJu/MMHh8PYZtP2OItjP7nX/vRVGEv4Q/WNz1sGi4nhvmV/G2lv/n3z
gfBxq3A322W6ww7cIXX2obLiDiPN0iG2RtabD6PmfRGwvRLiMecXAg2uT6i9eTFr
brd15Q1id3cijQltQt4Y3XXNSVkCQwpKaQA8zJgs8luit4A7G4Lb1uiU9e1A/k+A
rg+OrZCeDP+WaFCV3FQk1wUBqUumMiGzIF4nm6ZSARM=
`protect END_PROTECTED
