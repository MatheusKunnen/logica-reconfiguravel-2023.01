`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1IXM8KPBMctIE4ZK2AEy/k5wz85B/dWzx38WURq0lmI2XL0OE5L4StA5W7sfS1+1
uHlcEMnRhxqVTNlOQfz8IKRImy2y8JGKzL+mqdkIZ1oQnnE5iU7VU8FfoSMXKCZT
8t0qa/0x2HcnE6ewsaZD9uCiQVYqBrUM+2cSrsvV6FuWUOx2NEqPbkDE1FmZJAmR
+0tFfqUzZv+uhTDOfVSLIOUTWpklSpu2gp3xJUJZ9MrjoKAjXymnaV9ab4kPYyTX
dTmrRoGhtTwMw9Y2yZaJxSbiUCzD2Il+mdf3FJSZ8RqLxcAz+AVB7cQhQJkrVIVu
JNEWn3UQvE6eEHbtDE3/8Ux0io7jZiCSMt80Hqkgw1Hb33cKyipZAqw7IIuEijs7
iuVGDh4tw8Z4P5lOcbl6vOKtzUff5nSUt+7QtpQKqwCxllBd0uucfPzFIlXcOaO/
/g1dq63YeWL+oUraj/MV6HWS8Ea4Iw2usJYo0Yvjj3nyuIOqNPtnn2v/rhWBxkMY
vxurntJPvalftBOGkHQNm4l2TpcwJCcBLVQksKH5rdR0Ko7yZUPvKI1wncrsB43q
UfLPzB++ncfNpdJ4Tdb4YAAJLKrfXcV+ps4gPnB4J6hGEZditcknyKsEGD4mnWtZ
SN+hCngZQ/czz23q2uTg6+GV7+mOzx5fiP93qVwbamL1yWWMnIS9jhwgIEbPhXpW
1Lnu2KOAlOzVixLqPX/m3+HY0HvSx3k0RGdBcuE7RvmoO6gna9prnBOuxl3yY2rq
SYVOm3FnD0zmL+6F4B0uTY13sVBDzTAjVM7uq47F/SAlxZ3hfAvyHUrkLvD/QwcY
GEah09rSEWC2L7o3eGh36TAo1rmwVVZhJpxrzQA8NypcR//yxkTlE54Kau4n/LQo
RODuhVtmAvc/oT2x/o0XuHhZC22O884V4UC44zqHAUJMOxgQC8hG7QMbcXbhYJGq
kxeYcJKWOmN3i+ubxi1Qd6Io7AYyI2Mgsn3kY7DL6LJXZzraRCFzUgF373ueS0yv
bhQRN2VeAB7fPPm8iubz0xV6/zDh0+2txV2uut1Alf629wuaWOv3NEtmo4asLNal
xLsGuMOIMT+ivPSssd0i5cFG52ThII+KI8VZJwW7f7l3EJYhyJe5lOYQX6NC4Uo0
7Vx0Sv0BURTzFqBRamukWdjHAeixQPUzvkrmGjLH8qO7CnMtb/5TywUJwCBTmS6p
diu/iLXOEFUC4uHwMran2VkVqh5GYJX/Sn0isB8F5MD4qnJxrLsbi397MPCVFZ8z
Eqz+lxKFKQIDX88hM51cK4q7R2PZKBJgoybiI9JjkK/yuFq/B1HluolfP69xmkVK
XKwUh6AqupzVCsaYTweVczQQTDkUq1CrK9ojxXdx66iY9tXviOdZr/f3dGHjQnZ9
kofuP4Mz2kwozd3L7u12N1X5Iy2+9O2TxAw+63XbVS/6sdJIKPE8d8CyiIA8IM7H
9dT/UTwsM1afBEB3c6Mk9FeVnKBYJRcDXeJtD069tOOdNksEcgVTIJAyUdfZgGoh
ktzYumTzgN9OmqpbjyotL2bokhX76GAwOr5dNvy2H9taZl/4MeM6hDcHDUKFvhyt
YDUzczuGIstxj4Y9OY8HL/YBwfspOm+EummhJt0LW1BGqq91V7hJMIRNnaVb+O4L
bnPOUzVsycQEl/tWZw0+anxKhg/fL9Ptk/e3gBKo4Qch5QmzdK7f+3lMmnJpcdLJ
OfHgGk9x3BklbOGCuwWa1sm4/r6gRL8kC76FjpFcH+ckm1vpOlA3+Fwq6KjhRF6m
WSjWi4G0EljXedyrp4z0vSX9uPZv11ebLvhr1GRwCVPKG19v62qRiAmeqrkSASi9
v1pN0mlbjESIgVO3HIKwg49+kylypM2h7QF9VtYHO7Xt+2R2SmKVHpHEu/aTyjbP
vu4aHFVg3Gf6VsmGjEY1pIhQuMh3yCUvdr34hZA6kUHmImP+WQ8QHb8IKAl02IdG
QpmLjSal/xga0EQvEHOFhFFcrRIPFv5fMCkgJYhIBh0e1BtxbgAdET1cosKopSSS
9CJ+bG0pMWZ9TH7DC8MwPICEibr0sIfRYsMTwJDAAm5FlCllNg1+WmZcngpjOKHX
Ob2xQvQxQQYPojMBy/GTszMQCxA6zQ8hq10lRXKITNHqc+hE4lE3/Hw3R7jp/nRE
wj1VoPTqFugRZnGyN//NIVFQN1XX5YmdEzxqTK6yG623DVl9GRErgQNnDpyeVymQ
z76NazkONQP1X47E2DLH3r+TzFuMjZcJK8mOo0wCnYplnMdiMbXK7s4j0ZriSMB9
WpkVoYX+wt+XPIbNbLkELvZD2B/NP4o4WM6ENqZcuvfb4M39iMz+oQr2ySCvUtUc
O77U3lM33k14Q24NthHoJK8BtBt8XUA3xilLUXsWcF93i2wi7QqSomzn0t9lXyRH
iVDgEiaQZtpIqfkUhQAPa91hBVb27Zvxwx6dZNGVuhRGIfbkATNnbCW8ql4oHvXS
+dP19Tvn39PZTflTRtfBhZ5zFXPSagHr7ng/8u1mUaFmr0svY8TWbMc+Rrmc3Tjj
eS9cnEgMYJRKsFkhYvoT1ktI5+9Qk7vvI/JCTk6upHqvgjcB95AfsIAL0dCspWPF
mfG7ayMq9gNsPmUdGfXDtab8bM8WP2zU88rawsjTG8liO3lNuppnNRav7PZ+buZk
XC0T1pz7FMcRPwIOCLB/+iAIXub7z4g1/bbOkX3Sr+VSXpwC+3aYBb+Gs/klwuZk
gi5IihbJsrTbYsE8Mr8fQ75nkfZS7wyAMSfeYuTGemZ5Tm8pRqBw84XQ5uIMoSf+
aGUnWbnbtvbrutk/wIiaH19QsjfTdf7sNGwWy5pqEH+wUV/XLqKhjMKFvJH0CKTz
U9VjORL4h4MrqtMnJQlFcozUNOdnbA6HbMlBkIYDGO/kPYTDmpV+rtBN/d0TryYY
roOSY5OOkeyEmnSNVeowTIoycVk60ie5BtKzU+JQPDzhj+iy3piazGlCHXKotXbC
IEu4C297SiclQXzemujCSUAxzZozDfQUITS0yKSG7t9G7sx1aZfaHfpOXD5OcYBe
ffd+223EAtbYo/6NQQYT4TUegxytITw2z4YN2WnoblAEX4x+zlh1BTdzUq5vkN9C
3Z3YcV/GYN5wCYMnaiUcuOQLLSPeJDSjM3e8AhBiZbCzaFV5AtLZBNnElbk8RXgV
xuryGW2xaUmN96dO09yt87+AVe8mPhuXylqbFULI08ZF0Rqpmx9RhYtAE1+tBLnh
DHxvaen3NNFEo9Xhd8iVCrf5tDX4i6cX0D+HMAKiivEWK0In63K3t1Vs18h/kyE5
tBzgol03DzKeoo+K8cnRYLWDNUsX5GJHCsl3IxtEdouwwcvH+B1FzhcmSoqVe3li
OF/Z3vr4PvyGtRGWHdHlJZbfdQtn50Ow5IPMTklKf5Y/l3NsL+LEtyc75eu6K13u
hdyo27DwcI4PizkOL2Aug6zF5lVDPlaIr0QB1ftFnQHCPLQM3Bpen1N1xCm9EOXa
R1RgMxH3zWSINPxM5i/gDT1sqWxlLaQH059dwOReOmyvNNW/Hq1m/WiDumaKTKmS
gt2jXoRAcCh+K79gqApPSrePhUYGlCUaFS2j0cBljLrMAEWntrAzv2/ZK1xIxj+Z
7xIVxzMIGy75cph0TMW7t+YU+aBTA1MEeJzDVUJRptCzIEOQHzViLheiYKDWiJod
vXLuxLn9qH7QET8RdIk4IHyBrONlGvZX6sbpsixvnn8jJq0RGNlh9HVavi6Io3A0
u3c7w5PWw7YGyjDGrWXEQklvEQ+O1fsSw8jZhQBxKUS/1k2Rg3A6fOJo6b8B689P
8ybY1ziLdILWza2wuj/ne+ZmE4UViM4xfVxfOPk7MUGJnw7Uhls6VBNXJDFPuqlf
suu0Smph5NjHKXgQrWDHVIukNeV5ONvaeAKi7CT2V4azWGCA0uF6CGjs5RMWcaTX
jxn5RGR3AmN2U3B16eDk0s1ESK3RzGhjX9ZRdXd9JLF4RiNZy+uSQn68yYtbTAT9
kD735XDi3WxXoboWmrJM70HLoaiFBTZIkXYSZu6jl182bfOG6GPmAtXLnCfn7pKL
97FAnT7YBA2Fp23jvmoh1OBB0f6A5ltBvU5enOszTswizBgNillq6ofu2CV6INTF
AlHhBwEBHnNTf09sIl+WUhQjtwWCGhNW49/piWUne38UL0CfVSoy3+ZcXjkf0MoK
krK6ZgkxxQuNuBgksOy5gBghckf3CcqFD6mzYrlH7PcbKa5hwM6ExVgg+kFNqLe8
pp+yvXHhte6KpvSeXMpj61XcODT7TbztZAOUXPBig69DOu4B9DRO4c9SUUbotalp
r6QcXrBCl/EEJQCz0cU7iFTbPEvlQRU5gds4nAoxGUtmN8S+icdY76KlGEyTNi/P
CC9rjSchTk9xMptzx21jGEamaiNoWwU49tLd3lCaR4hSJKIc4yG7tX0rUM21BWOO
GYI0Ro76cxIg34bS/ZrIekp+UCgezFY3igUXztI6SxMGtVL7/PcvIG5Q81ALv2c/
M7vNi/2qubLEZJgrPp8fxZtuwXbmpI3HhXC7MIql2HWsysGtvL7Xff4RUV7CwjMj
DPdTsLh8KIbWk64dFbBiVO9OT/oBQxEOYb+KVgr7KiC18kgzNE+2ymQFmnfJ+aA7
ZjiXU53vAa5jI70O059WD0yD6vsSrQjtIExsdrKHpRJwgcmJhueAng0TF0uRVHkt
qAoI+OXwN9r4GnO/mRTnuQmlifWVVBkzmvUbGS/vFqkLOEQAGu2ITzVMpG8ZC8g5
440l/K6DpW8WvX43Xg80y/0YfKI1r3wPCoTq9oe3gtERGrzZzxbEc+6smyaUo/4I
cZy3I/dmMQ3EQNZqIOgPSwb5Nm6o6tCFmSiaKAMD+wDtQiDDh1HKMF1SBCrVfXhr
UU62qz5E3rFl67izQ9Sabwbvuf2ae6YGrhNPnVvyZY8S3cHKL9H/Ov3XEm44WRjL
G3EDz34Tk7wSCCtTMA7MltfX8llpv2o5ZvMheppKWOYIHo/qCRCK/5RfZSKK2C01
TAKHLofBt4wvwTIzyRyVVkDwmIiuO6uePNfKytcxj0poCAzzeSuiKc5fsWE3mVCl
Y6BCv73iFtyBWkV5MphLDI2bszx1PLOBcP/PvPp53AbggjJHbX3ZCwcy9Cdbx89t
OFEqBWgWjKDaT9oHTvwZ4/TWDSIonVtwvGrBn6HV64OE73iRj5jql5Acn7ogyy1M
tWP3AfNL2LGRwo+Of9SwaoQDLgk+qq3LKLMtNcSmu0ewyZkxl97nakXJ4+SN2HIe
bhMn+BquteorjywOybg4s1jpDQOCRVB2KIq8jHMRoq8Xivsfa2vex+q83J9JYYPo
YcmVyfSeL1L8HajczELDHJG7lf66/upHBTtFSlFtYNTm9D7Q1bxtRpGs1+zfjVjc
Zn+9Q68H9WEpQxiKKIEMYRQJ0TvXGQpRHxTNC/b8tymmAoz9iMRbxJfDRyKPHrwG
JS6U8K3Y7ltj1+JdP8UpfgCaGbFHGaUTUwBktXOAD5edBM+R7rAQJVfBg0Qtyp+B
+/GSm0if55ZTtmXznxSXa+vU3/jjSBtLLwIiew4zNFvHylGd+BI2VRJC9k6xZOn5
BdwtjIk+hzgumrS+s83SbYa3hDgOz6npGwrLD1QxRC7Ff4sx23/XHnuqfkzYZohX
`protect END_PROTECTED
