`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UTi5LQB/7cgwkb5Ly/vn9i2wnPoPWIPkiw2V1bcymu+0jfilVCt/l4tMIhsUoX78
TbuFJ+XujbtsHSbrz/z5PUQaDRCX+ZqYYoVY2bR52JEMoOB53x4ptImwUtVCNTmh
NDYecH8dl7uC7WWsRPTZ5xxoTltNl2cPn/AvZVimf4IdisCAWf8Lgn1R9w0ijnWZ
xBF28Q90+vsYiRxjSro3ISqs90xasNaDOWEq8Me1Ie6EEZ9PvOnslN81L1AB2wkA
t/0QGg/tWWy6GlXf0/F2KexGgzZgQLMRoS03d8RmQ0/28CUayykE4nrK8cONvQQo
Rex7zXNkE8neS9tTCPv/owKcViXrfu54C8KE0OI1iYSfsWazA0IDFKzCNhCXvp5f
K5p1bqX4nMA/5S1EGjz1N7gIQ1qw98CnCfPAUvcZVLhqL2MIBLpJa8z6mlsB3J5z
suW6ipQgM7GtI3o0ebI+mlHlwOjOPNkXMYPd+yWz9GQfY6SnWjNYfQdhUnFkPO9s
u36iuoVD4UXoJ5XiJ45h72ClFMLGjh2mYvOx7ahFmSzQA0xWGdYfgW1VkIslIo0Z
1p8UXyDJkzwMPWAuwyHv/6XE/U6oroHIbgzHN330/Gv0kETcPweNBN7syD3/KTO4
Ubnk38klYf0+IoJyIWlDyWnzMFxsBUnc9+0Ch5qqXtrzthvZCe2ej+LC+b8pc/LB
c4bBcPzcUF0GbFYpW23vzQ5WAwfNvYlQl+K+R8sgebPSFag/reYreAOg3cCGAVpy
LjoHKYBg+C2rXUK+nA2780TiZW9XWXiPiL5ro3gTlksCG5G0bsI2JMmVVVFujoBM
D7TFQFTOQt7Dyh7y++1dDwZ8USLUyXKqcrUKkaNoS6mgb4z1RXs4B0rDN+0+qEeL
EcFa0twyF77eewOaP7Cvg5JMBXkFhWQDg1LNbLbSJdzauzZ9h1bRu3bRMuE5cEF+
H6eGkVNmuBRHeCss7q5gfyp8wpG53cOkeE50mTr0bAxNKGM0aH7jd8Iq7AvCwPla
wzpG6sbsqQCo/9Rxn/KkXP8aJT6Ixlb3Y+VwBLDkSoAKLpWGooom6Wny+BqgYvau
abSjVsLjNHuZyBzTZ0KNWmLSJFkV4WcFcH32WoGUZW1RWZBxfJD8PCAsdK8aTIvg
S5qQ5UPW2VOZqccYqxilzRPPRM89jlqk3E80zBxAH/tw+A+WByVVS54yh7MC5iqK
9giAEIp+Rg4PWT8r5tq6muKVMGapq6BkSXTinUV/9yW4rqPGTNtbbuDKqofWrr+j
XJds/H6g0xVpgu2QYT1hvPcKXmPR8tffqHx0xwWMIa3RdiucEwyhF9DtLi6z+6Sa
6mtJYmqGzzWPnGY8bsKn2fC627f6INrePiBE99NhDEv7p3gL7HcCKyHApsDmWK+v
JQopKgvPtBynLqdy+as35H1LQThq1AQBlEAGzSq8159nKKFNu9YiEexcYKpaOA4z
AMR/9K0yn75/iK+mQ353N2lvy15FNPom3H64P6+JsaqHgDqmVykycmRQhCpd+fhm
NCSv5FO6gFoaTTJTrOxcGf1AuBSKHPkN/gcbOyu2NCV3Z2rEOVtgX38CKX1B+i12
tL7CA+gmIszdP/TZSMXGK+p17rJQ76Ayy+gCtdwYToe+viNq9lAwKwRVQ4iKK70H
tnG4qxDuTz3nPsN87pbB35UW8TBLhtKErTE91gT7tgB1tffyRBwGNN2YFTVeBb8q
29m2oBtBJnx4DUs71lhZcnfHBGcv8axP8fI/MSlDuuIfTWJdonXODJVF7kc21dOJ
C/LNq8PNsYB2xrJ4V9FmzndlFoEr1VDrse4qprnhKMCt6fqFRUj6hRY4yq5oT2BC
vx4L+UKtHssGzFcOe7dHzYEDjvM4iubGAVW78filFPCmC70xdeQURw1coVkqLD+a
4zdzhJJT1V4f2U8fx0oB4GHErw/5w0pm3H1eNYEswTHtphQrCXWs9v14wUJyH0Km
PcerN2XyS78ZC4o3zxBCyb+rXwQClbjkc9Nd4dcpvuQr7WFx95UJGib2MHm8QQz9
ZueYnuu5YUSszt12V6IAlhhfkC3dMBl2hESJoTBjqV3WGFTipWdSQb2DUnJkQ9rG
ShtYYtO3cPEtSl2RxzcK5CFBm7BxHZESYc4ppExsA0JrL22KHQ4nmsYz58HvvxtP
QXrYMAWmvxeyt1pQpY76fM3QFCieOOmEz5uieczhppkx86HsFuSQD97C2Sa6H5pC
nfN3ONbpOs7lgLjuSNzSHXBSMfraOR2hqaqWBWy2fk+Y5pvAEuHdWt2XnE1zFJyD
hFEABEws50B0aCPS4tBkhpxb1NrA44SMeMJ5vak2myCYhc9z8d8bT0mN9LfVaYhW
n0NAxpbICQZdYWR9HmA6yEamVo6DlOozF9ELp6xUkD24PE+sencaBpH1cddNXKO4
o7pJGt+k1crQLKWrVdksyJWix8Ct2lt54QbGYek1+fEJlwfOLVEkwqkfXt+jo5UW
B0uRD5zphIVdqQF1XHiaSJ/RCXIGy0RPdyOKcNy7t2Lkm6qKAZwjTo0d9+vlaeLg
Tq4xAYoTepAWikJp/7vGrfc/HyOUQEZmU3KzHX6hzewX0adzfPwIKfp+IFUFJjSp
yCQ42bc5HSwkiWgiikbi4x5kutqXqAYjlfKqwJxA8i0M4bXG/Cum5b8OKOnb9LRF
k+iWK0/NX2trWyk8/lTLjkt9VR5nTQDmOfJVlFuqEXgaXIUnjsrcOHdRIEz1fx4l
PWhUT0BDSJTMxRS9Qz+Ova1dsLOozFNqZWNxrAiqrpNyP/hKhoQQ4DZR+kKgOffg
rY0SpR+5zmpwuZiHIYsAgbDuNhVYzuoqnZLMMXst4YNyeN4tJeFd7blSWqfuS+HU
7zXBbI1Kt03BJrkYF3Z+KjGPQw1zbhdoaI+VLK7gNVY4L5GSGYL8Hp+LiddRYZ7y
psj4rBaA+WbhuV++vav4DzrQZi5UqOyp8/mAbpT4Qot0xmlI1p8QfP0br2I8Ur/q
vMKW0bYSZ+Wg2J97UXyDGKbGnpc8W9qgldIL4tDdbdR/UPunTJ6d4nkPwxJROJ0q
eP2JdIt8RuEsLQ3VaGNbVkInHh4eTVSlZ37KcOVUTQrGsMGz68sKIdorxCd6I/fb
b42bt5EjB2aFurftCm9Ufib0e67xYimA+5edttTVAZarZkjworI6O0cQwtKJDZRX
X70TRcI/iRtUazIPRJVljaAd8AUPHT8r60H3ZhBo+zumOTHb+IfQM59+mTwbnY1X
+HeFdHNQoQ8JIPWhItz/QpBYpauuzU6Whs22AsiYpu1czU2YNO5cqJFHUvrj8ppT
2aSBOTWJM821/yk9x5lJoga8B2hV4eH39AhEHbEkwRPRWRgXLi5tGB5aTyO9fjVL
az9D+7BooGFYaxGh+71xKfEGr4Z4sUXNNDc7zOdv2ntLOXQudXHH7xFkvbzeOzf9
JlhsUJzR+zaGRF8OztTm/RLZNlKRR5s6735JqvLsvfcF+qSTimsh4YiHNj8M24bt
EsB6WtOOs0O1qsUBIqMfTy9EhlT+MyTBG9S323+c+s6RC1+8nuPY5UMx+gJbRzbk
h3D0Jv2YZVKbo4ZNe+sZCInhZZRADCKgqvnhUHsO1CKSt7uez5invbKN0Ltgd5MH
RmGzlAOgGT31/tb7uJQgdss11nnO0eOlc+kEOtmXgRWTKHJPbsZWnv0hnDf9gwjI
oyle4Y9s/AcB2FAlKWcsj/8XXRgHeUtyUQ2V8y26Zhr712L9quCG29TCVWJ+1j5w
Dvfk5pFegVh0V+pCZi770alhX78kpYyJ7wEjVcyZqbqRNGMLXwV9OQi4XIrDUFsc
tZ+5fvBO3KPRYsCKbJKCdhbmCZ2+fEyvXMYrjDTS2xo1awP5J2AIF/lW1XEJl5Kx
XhOuGSpbHnev+tYfFEALf/GhgQ7bByNCi6GGUUykCVimEFwE4dPjX9/+R8oHtt0B
FGi7b3Fdgb0ZQ/M+1d2vtbjSeuFC6BmWLdj2sPi47OyRlfC30NpUESVxz18l/3kb
HHuhWC7mJcZCsuiL3QcD2MljJ902Na0pKKInuixqUbInFYp4cMIQ4KrXBjGWa3An
RlAuaut2yurVVHBYtD7mui/r6/ck51/XOg+p6HYSYZDawUXnp7/NHWhCoZWvVezu
s4zLXkggfhEqcksYOrQ4CEVKBVHQ7PSMd3Zlncci//KvGOomSjhMT9VWCyHNoDMb
4syFSy3YYDqNUFpRyHbpl/VwkCtZN1J5YrKnoGo3cNwctSJYMA2KJ95XaytfUw2e
dZMUb9ieozcidYgoPNAIUyGxo30MQ4yKNgvDQr9bOzJ5s+dx135dARHHEOf6KUvh
jiVln/iQIElRnyKUPAabcQCtuH1eROmQ7HaXnSY/3j6hhGXM+aObOhr/GMZfOX29
87xsJyDj93iWZn6IKlx6MnLPoXmcyf0eo8kELW94GmjyCnA8bkZLy57ro+E1RdPA
P9g8R7TIMPSOB2ehy/SGrTm0PR4KD5pZ06WLrbmGFYnIf/RTC7lFtBwo2n0jK9Yw
fYcD99VfAYhJ46w9OyhGZDLoN6+Oal7+zhlL/l7fFamSgwEWPnQxC25q4ONa8UMd
bd83OvIrP0vJWCqC4JWE1qMPkXj/zCiF3kXHFoUq2Vur874jyo+T/y/NKWsWAXHk
sQKVon5BnKwScSZye5lnIVrjfAloMB5ZAeqpkiOBrhSMCehE6ApMD0ioSvPmV4Jq
I0eLX6ekqFHmmHN8/a9mxQsx96ZgWU53JF3JZ/y0LMSspqqO8M3hmEag/TSuItlc
v3vevSt5ZGUjt4k9scRneAebbbWA0FL5w7TBwogidrmLRtaJeWzKyZk/SHOJOcx/
BzpwoSSUFSMpB1Kvg9UaxJS618CPt/YzX5i8ELT5f4xu/i+QesZIcm1u+yena9z0
Ic7U/cYZCH3gCUPdADTINk5+WRwLrhYhRAdqJA1kampQD7eZZw6fK//sp2R04Uue
pZdMtgvstalIJTnYW6b5gIvS4nNV0qQ6Lf6Q8TMiNZfYLG+9MrOFJ0Od7iCobPXS
AQ4zVIcCk8acN6IKXNSYazJ2FWNiKD5Op+ulPSA9rc2HHpEBoWsu+VMpEWQ6VMOm
Dytxgflcs8VOE4o8n7mjtYRYC1ch94fbUEOiLvpfYKnSK0lswjlQV0cCCmt+7vOl
ZJs8YWNpfHTmXZdIpaWSeYbuUrDU8Yg7CzsPyzLliOvy3TmPirR6yXPBJ21J1K9D
04HvXL5x57u29UdJlgCj17We2yDvLFzGDKIOnhrsGWQuu7QlmKuCM+2Wgi+09ek4
uL51tpEJ36JA6vr6IgxdKOJz12tXUNAOruHVEKqTpP3E5EZM/x/HVAk0AajkTi3W
hAAhz8kNavuQseJykffkAyLjLz4ijrBulGTHEt/zlAq44ceVxNtLFnwbfznBQTkU
tSwAfV0x9gkZEEleqoj6LbFk8JH1LcJXXWN1FXJmM3inazp+wnIyZIExUPNcByDq
B9q4RwUP07zjHe5n15mw7w==
`protect END_PROTECTED
