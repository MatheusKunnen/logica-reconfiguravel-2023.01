`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DaBHBFHF/Tqd5Gw/kg0tFQFlrtnoLO3GAiH0y9SwQlth/cT5LGnY7MkBWFiOmDR1
8je0NreacIkJRzFQRD0I3DUwVdPsKM1JsH8SeenXxhDAQ5Bpl0eqvj5+wR+JL/yG
qZSinbI7QL8FmossWum8wTZS/NFPcYepSPy0b/dtKJD0SFh/gQIMpVXb8nLF1qTK
1LCuM4riFul2jrGu38GsWFdS2+6Ww1EnY8QzIsn2xscOEo5ogkgHZ0oz1dFebbKL
eApLoXExjbQgn5F0WhuQlwmGe0E2k/rWdXclVFH92w6abZpy0t4NlXQ7xgHGJPIN
Dlce3IZQwqFd2qZGi7TtVLltpxc/3V+iMshCnB7uzQ3AH2LUanyEHeBigcTDvPas
VXK5Y1VczAHhyOV4SEAmnFqO4Afaf2jg8wUZR4sfo9FTgixfhRvCjXCN0uzIKKWp
VzevZPIc61/Kn3JB4zLxmgrZlin5G/URJVshtWfkr6oQyruUhQf4Urrkb41/8aQJ
KeQv2QaQzdOSvfCJvU4Vtoo2AvCD5BEQBfeaPquUkmUEdw7XvfZ48TfH2UvVMX3f
VCyTULlqT8kgKxnwGgXMkX+hiR9Km5DPWhET3OqafjY=
`protect END_PROTECTED
