`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/SvfMhHeBWQk9uUD2IZ0O/AOEA7plyB9GHk/k18C5NunrKdqo1rE9Gmyn9VvWPM1
J4M6rHCHKOiVX1k+z6CkmmaNRDUub+962FsiCL7rFI0eqkPOk5sGkvEDgI53Xhzv
TW+rqNiOBPJipF6zhzATBBuwad9qe+byaO6GWwJ8dHQHPDxsWBdExpzo1foNYSnt
89BnfGZ6Nk3N9XRy4iNSZNVEYfUQsQYHJncunU4s4QHGG/vTKhFSVSabXp043XJp
+/nXE2FeO7RjAUewFlqP8wNdgcRGA4K+0WrjTcsR766MmIZ5seDEVFehjMn9Bn5m
4hFfrOqJ9dvSBdj8V+zgh/aId+FLQgCYrouApnnEqIuYUYKPox8sBnguilz8FdfT
pHGZIgNtzSVN7f6Wcikonspn8N7VtyU1Y84K2bXtnwzZyQz26BNOgDSBVSae7RCV
aWycYtWMzLPRciUTi0ZxJGyT1SxYPz1G0SRnv85EGGdhxqXo7zuTqeeRv5Xdm17o
v3B44VuRd0dhAFo+3+YZEOMZgYiWQmCle7dLhV6YzM7HPmXIZuoAcS42kfyaZpnj
p89nYUTer7rSq/3dq9H+nKm6/Rc1UFe3J8dL2JM20LKK+aHd2bW/9JpKlJUMPgfn
XIdE78asf7XecEUl3DzOdjR5BeAzAELVsbl9gHKnqC7gqUWYO9qxROy6RnpaEItB
NPLsfTI1iTlwSkClvnlP8kVnt1e6L2tSKoTBdAenT2GofaPoxzkEfgWy2fNZD8vy
QVpIq1P5X+8zeziv97br3B9qxI5P3FK+yjZHoECHFHOfnSFBkeElm8TujVIn5YFS
Fe9yS3cvwtf3TQl7C1F5zJyZaQMOkzyiWlMBBOHvavXO2Wy5s90FBfbkO3zRXwbw
GSz10agDbuUck9iRVTwgaWKiZm1xSfLTtWYZ8fRqs6nZU8iHDN7lj8OzzO4LQwWv
AjiZdohTm+AzupwyDIdl8JkGGH+cbV6bN62xnyE2XENG9slMf3lz+UG8fF9zECFD
P7Cv3MEBC+GyMplS8nRI93ktm1bAsoCNkxkuaQmvhb25Js6EXgdiUuvMgxhxJ3Gl
iG14DHMGJExLaiAVhifgH8DKOJtHNjf6Cqy8xCTBxLGGuEXZP/9LHhFPOoDzn0Jb
qPPd9sXMH3HaKec3o9KjglcP5JDTGA1aJ4OEbCSIPr5NaKwEPgoj5UU7URoVAIv+
ofk2LzmPHNaN7Inma/48oAz0ePRutOoJYPHw9nTa02RkvPLd+D+Qln3uGKKDOMjH
znt9IW94CihhNLQesCxRJaejMCsYJYZ0NgVbcrNRF2SErQbMLt6UCJgcbib+6gdA
sWzurv713mCse1aZYvp5CtHBrZcHQOH5CLzacvY2wfnRTfEqOLs8xjiJIj/Jd8r/
F5RZdjiG7Hq0Fh883XqAIDlZl0KIjldrBQ42+KD6/nusiu8aYmqXpfGl+Ml++Y7r
8nRq2ehazKFWkAbRHSI9zrs6iE9+m+6BtQWB2hocDbbtlcZfce+6/dc2V43fTJCu
/7/2uHyN7EWoyPnk9KGouAstcas43hW2d9PVa8U4sWbAIVW5K6YVNpF6YtRxDsPD
5fXCtBDXZrG2syGcavLKKaMUovfXplEY+Ht1/M8NjnMTJ8FdSVoAyX+hobPXyxnR
srWgFVGRPaSyOsWd+brBq6AmCXwN8YNL+CWqg425WU3A7eVoSfVG+gwNkK/qwWKM
SzmAJn5Z3BTv6+zrnBkCIsNOeQfFC2GWbhNNxIZV3tWOznQfe+XR4xyTDOJOlIiL
KebL0Ng/3ZWYkf/6joeTBmPyq7Cf6D+AX0nOTzn79H8tSmfGHrcpY2pCDzcxShUF
j9zvm5IOf80J1VrJYxkPWg854jR3qXjxrdM/ehV3vpp5lhXDbL4/VZjUHEX0as7R
0YYyPexDXQlKa0nGS/SvT+E1n6kB+3bpxb7KKig0i4pMm88Kl23wtRnUr6BCHShE
uP1xSMzjLHDPLBJgJ3clByM/iljYwxKsfVtuLr1nV6fRv/1B1B+Us6mZx307O8ow
Io6vw1Dadpe4e4T1USuk+CoM+ao1yxz6Xgv56WGs6DvnT+e4G5mpYG+q94Sibhmb
vHI954no72mo9BF0jvevts1I3T4vAnaF4uCYRVedIrR3zXWJysCySSsXarBUhDFk
0CzxmRNGQfmwFmHKjsK4gPO81VxUoDWU8eybOUUZNmP62skvMGWXwvtnhMIlYaXL
ZE50MsOIBHQt7vTKmQREMw==
`protect END_PROTECTED
