`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HmZKg+Kyh1vvP+lz7W+uZscHyxd5kRaQtjalgATNKwMWfbTJhyrN/5KrXJTOvJh0
d9CemOaVIa0SWy4+qsiVBomy5/FMT214R6WVtJ3iER9OVtxn7sCF3AvecNLqXUUC
mKtFFlT8upIjRv0d9xPDR+45yi27aKewg5FTVuSfMsxgu2bNUoJqpP0YdOuxv0Tx
DeIKsSXOiaKEWSiw4JiQaGrXmJu2PKVrLVhYGtMfyMQqsS25fCSCAsehMs/GBbBR
mdj63xxA5AcOd3LOBdJSVVek0sUwBhfx75U2WNb3nLfJJHGviObjLk8iMnnoBO36
tbm68j/g80pF8istha6WjAgdKN8jIQtB3S5K/hDdI6oEUA5Ol9FdZVUZ+UPhgdyQ
0tdPrJGjI4AAguTd5n/XOFtC04/u7QT6wNUhsEAwu26eo8SAGgYHCtDToWXffM3T
WJcfmFPdvavTmDWzhzM5DNNKySsVncSjBWWfbohqudequVQtSz4EOnKYhSMUZgrE
7vczQXpKuPmw/nBS/P1bFKrtTunlajrJkMyxSqFGiByobxZvoFhItW22WOgUBbDU
Emo5wpVVPJahsMIHc1aoDU9iUQ5qRBSGwy8TbeDwdHoQ7f84f+IRi26MnfjW2R6+
UOjiL8xcwdHiE7svIyyzva4iznXwKbXA7Zcf4YhZKcULohuPK4uZ+cZYJRuJp+GS
/RGM3jhxQO6crX+pJxkun6nfoByskXcaKN/D0TdDR9W8oWFpx5iFdJKkKN8U/1FR
Hawy+5JcaLf2wbz3R4gh544/7/WYaRc3LkUSKWKCaXGTGlkip8GEvcmS975YA1+r
puiRkjPaN8YhbqHts/emzoXQIjfNKWZUx8AQsgoXCSVXZncOhn4NxL9rvJk1VII7
wgmnnfzQAUab0MiLs59Tc9hP6pTGBu6Nqainm3/cvUNuWl+/eKvrd+8DbSngq1MI
oTLZb3rOCqhy/Vnsqd7o4X/eTSmHr8MCcHC1tc4aXbFLZDuTiC4LgdxLBL0jz6NS
0oq2t72pEyL2zCBIF51YhllJ1jPnifviuTc7QbQiNqrMLYTEGDy38bZ5U4HogPfK
fKw7+bUpnaOUHZ63lo1AhKp4LFNumUwZOgMm10cYk7IDmnzn74wgMJl/BASKfiPa
2poxpdLTYVoK0uPVOJl5jtrGI/SgUKmYlsizB3WrzanlshCXrFPSo//jRNHwMZI8
dxUS6O/DeuazbTWLfBXYHRTSBXq4jVkBKS4dRO4Yzb6/tw677hRBveb4LWfhpzaT
RyAkvc9DZfftg3xQkfSrkCNaqc8TMvWvmn78NW4kZXSd5JQ3j38w48uaVAzT4pl8
+gvq+5EgXTYDV5h+rLHk4JK9HucWas7SBEiofd2lc/PQk1k6+/OnpMBI41qdoB7I
88MjlPUy5pxRNBvcaZpjLq1KIFQIQ9fGQzZI6nPFx0SbnUFZW0KlWR4TjwDaacUj
KgQrgzyrvTxApPVaczjfXSy+VEIPsGANyR1bmu0NfTxia6DUZM/MBmJx+gU97Z1L
82zeyphxp2SVla3o9hiMOdWVhME1Fv9V5608RuFXkpGrSN9BagWIqa20tn107oMK
rpqgIsI0x1gX5WfHw7isyhf8JqUaTSdGO9ISwbwk+f1VRRVzYiyKruFqoSsxoEiZ
kIUq2PjLYtyiCypD8Qx3RERBR2Xfy/qL32hA1IuGKXsXKB2EsO6ZUqwH5Cpc4bYb
K+SpHADCQRIbr5z6gry4GNUlYp9obmFOiB3AXGmjhgVieZh1UnqLIjnPAL87QpmF
XKIcNKu1BaxGX1EJj3oIpHmM1GUuDtOo44PebPkWQAzoZhuF9UyfmMcqLhWE4v6n
/7pz1XYufGrabE4LEqMY3uO1iYLtzRCLXJ7U9e39ecOtpvnoa3VlmfjPOG8ysjgC
2RItOnrR0ks5IB5fPann6IDiwsvrl5vg6opiP+ObJ+S2Z7YeOYv7ZqVdFSKrIdjw
k6sjsU1ZgBajo7Sjffn6BW/8jJoK78m6JlAkEmnT71D4ORpePQg5+lpuYM0mJl5Y
Ge0VsM1KFlGVUoJ4g9EJcqfinZ1wwEZ3FT4s3ugOMPO7/plsJegNMz67Ogi9rja0
lfCs0B+9J1EPvO5G7rxxdR31/MOi3uDiQGtriaTIOXk9EtK7P6joSzRRW7jfJi5s
P/IF1KReR2qTy6E7VELCYT9W6CNFCB8RqUo8OKGaWv6hgvw6jkFw/7aW+yApuWH4
xkheULPuH4Blgt0Q6FzMLpN9+FSCT3+rEuAPl0uzif933OEctyox6ocikCcHLN/a
Fys29/joDakENtEiuELop+NeBsiFU+IX+EVN/ayXssttozJYLLzpgandCQ1qW99W
RS7vxBAM1KZ56gv5LmxkCDOv6nJg8av9ZX8SbdxlD1AhrdiECU4eR1woQ+ZyP7wA
E2VhqVfSDqWjoAXKTf3YPPswN/LY03BUgDHsDXK5d8u6hbI3vyA07oCVvS9e46i4
+9VxNQjV+l6VPTywr/Vs+TCP0dIUrY0UM/1e6snkGS5ZZLryglYdexSSjRdCXhow
PfqRY7N0m1D+Fktb6HsKdVLe6FA/bsfBEK1XbVQC6BaW4QiJr+TcjJfBC0Zqb94Q
hs686zAlkxULyY3CDqokB7dlA6a/JNkPE7UsKb9aSnoKJneP2Y4+jHZTpvyv98pF
/qELovCyfSNxOcaJ1NZm3yrvobQ+k3L6jkz+F/nv/VnqftwQ3vwVjdP2EurkjJyg
M64wxQ3e6wEM1DS3tzCpX2KeXzl2M3v4Sgv+RTqbGo6tYLeUK/t+r3L3rHWjSBF9
jdqUBpslQBLB4M8iJtyxGhn0Vn5rP9XpI3WK+tv/qsaeepJd5n5IWfbozCI6VdwJ
dJJC+wm/Sm4MIjiQyCeE5LoZ7lpc86hLeLveCvEEGePGX7l7Se7GYfFX9JDilXQN
vnp1VzO0wZzUuRf7R3l7H9jb056a9KF2a2HXbV/4MvUr1T+u/tQlqbZ9345f2mEF
sGoxbcPzOjbRU46JVNONhtkhDLbGFgiCuPxzOXiqP0Q9V2/UUnrLYGV5uqmjDqqq
oPu1Log4FB7Ol+QA3plPV6TmWpdDh5m826bbo8W+OyEyf0wf1jcnspoYKCsJWTjF
hneZSa28kv6Ew6viNQYF6oRm5/+uxP4ox7qxbeeU/3NTfO6AxKlJf2+D++vsYHyG
Y0GWWj8X6zV4EKOdjX3aWtjMKvS/VzDNfPbL8wPaocJLh5Rtn5VNZxPLg4rcUY8S
gjGF7bECU5JVMQtq/pftyLrMaWHWq0RFMw+WKrGoVm16DLatpWRY2CCo7BCyyEGW
XAymEI7GvxT01EQObCIbUCFtaRNHh5eXnK9xNl7ry+WvsrGz1rrEYZALTUtO239Z
z2aHP1WsdUh8nLqUeJa1ZZEH1KV9zTNL5FoYzAKiXVGL9N5zXVsIpZOEcHiPwLFP
/QL0vcn5GC578PjT+hVuj4C2UR3YSHcN0qceFx7a5VxJhIP762AAdxCi5KgCHBGO
xdy+KuDjjoipZTI4pmzwWr6Kx7jndfIpI35KnUZ90vQ8oqom11q4iXsNs8+JHVd0
vIRiV/hKGueH+cr6m9NVkcYZBQdgyCfMcfOI9SdHbUHwxH/Pq18lpokav7c6f42F
6fJkjlqJjuvtLVnP+9xzPZHA1qoiVxHmurmIbJAnbUnQiXeUUDvIeMPA2SQ6sEKt
cfBdgRKO1o1L0CRzYKFPD7L5Grs7AxLrOYPbS6G8xakhN4bor1RBPtTxSPiYEJnH
oZkdT/Wb4tKzNJddESjeOjEtSrG0aGm+Dx5cv3xf0njZ9zvowFBOP0VjsGPfFGoD
T2Zxhp7TqnVF9rb0x6ZJkjIBZiBClUhKNBcGlVuebfpnARJmbDsRbyUXy9edC/EQ
T7qp1fnAdjRHtN3oVUQzcBAX6eXIW7BRV5bX/R85ZPhtcf410sDR/72kal34HNBb
jG6mD2HJ2xf7GIPKC85e88f05RekSisDi/42LVeLLK45klhDhe1cMjvTYi9I+w1O
IJKvoy8+jisvs1E/NcptrSVzXKsLzprgmimXGz621EKyeUc1g6FvSUy4iz3QXq1j
uom4hdwTUQjqh5fka4GklMH/xSrOKz1CmgXdhl5A3KmchXIHlVfxD4rbvPXPwgAJ
7D/V1cRu3YsRQuyF9SjgDuYv6cBoP4bH5uKF6rkKQs1j7KrdT8dN6B8Ro8yPquh1
8PfG+MGQqqirspWkpDA8kO6z8E3Mw/xQhAk+NeXhEgXr2Rn0DdfOQ3hYNtnQvmZh
9xI7TFVvKMTvVen59OyVxdXybutY3JPCsh4kTWPG7EFmbTGYpyanBiFQ0HKBTXu5
3LsOgX6dtu4W6MDUyPUtt7aMK/opT5N2vqPlm2OyThE6FleRj99T5SZjYdfTH4wt
FyMGhIdIhBY7ywKiNIzBYbu+zls2qsGUHEg/lvC0Q6+2mVq8yAvAPc0x5q2lp7GM
ERKrPDMCiSLGqhOWCYDVfgj9GEz+pebjBJR+M0ZGiOi0urkRk5M0yV+5o//dvU13
9SJSXOgpjvZx36e3Uq6WG7XxnXEr3Ua7eGrvmklg4CuFAqhNBeMpxCXrGytL4Je2
8l22XJQ/TiUKRZtnxlfFnQY/Zd2v5rbWRZy+p5c9IviDCc5t4/A7fEd594H/mCYZ
2E1hduaIhxWAD2+6txikUt6vVagPI7YVnibpAbHah04FktA7lHCJ/79om1dfcDm9
xKx7d5JOZS/PuTGrwNQbnJfVA/6GroNds56rhUwabPw86gxkKjB3XuYyRPsgGvbk
11Fdldk4RiqapMz4Dl5rbK09Vd/12AvHl1x8ctI0gPsL81gl6D5liHb9Rlyo/Xrm
Nt4tsaYBid3IC5mDqp0MZz5eZ2wSm+/fFQe98mUbI72c0w8C/M/x36NuUEHnzUUg
ezfY2zJd1QWLITWP87I8DT9egC+jUNJ6im9IpSs115bO90Y1G2in1C3QA8zGi3k8
61zmnP2pW9OcuiZSTTschaGrs3ab3Rmks019tDVy8sRSYUTfsQwfnxp7pY81V7CB
kTes+ZBVVcDcwVdEftJV4BEFc6qisdpsq/lSQnYTQGVG4psDlWoZUOfcXHOwgEvo
P9DNEiJeHD7n5LokrRekfZPDC2aAd3XcnFxkMYy8rTFnVFSw4DFC5doZ84xXGXIw
XDxW9XK3/GIIG/ZzBngGtmMi0wmXFNX2QypUoi9w1zkROTQs2KSWzd28ASx2zmrh
TZPOm0J/rC4gtUtQZuK4J+pVhZIxZADp77cPnBQJumkjWht9Ab0pJxRCPYAh65vS
4YCjPVVp4xS8zEJrL2nk9asAnDJzi1TY37AwfAtUvxZ7oqiCjWyI1dePytMl+Fd/
eNhUXiAYyNKNwjAnzSBvs5FFjosnI4yX7FV4pxQoeE2U7tyzPv7qi470XLt/xXUP
UqIdsHULZdF6Cl5xsV1A9MVlfZiaRNoXxfFB0993pASGxU4M0KXubfX+uhhoJsid
5RvS/i8M1Hcs4AzsSSKI/Ngbj3FfWM0DxiuNGC8/KYD0KGGUzPzT1iy/095Azsti
sPxZ+LGh3NqEtBhxjuRTTMpQqgARxadJLvhkh8NgjOlmG3nhO5fPnaY+JxBq2bUC
lsQi2qtok/bsfJoujT2COXAsq5jmsGdm+8ML9fnHEk+NlES+4olQtfD3r5xbYmET
PrmqMGWVFGhiypC1GnMmUQEGr6J87g/+YAQfzi5EJCTUwR0GbJU3FOF43HK/6iSC
bX9Ojom0rZQRR7nJi2JdyBKhV4qYo3sOn3T2ttiU+M/WPCpY8uRuG9aAMkpitryI
hHbfoCZ4XzUbe0187dPYViBLyJ/DXYvfLU5HakOZ03wTH8WXagBSNZN2q1LVO1Ae
Euiu3HUH2JGuIAvzylzKJoR9u7I0dPdGz7HIy5v75HmpH/7RHXffRl+4VGIVSr6d
Ot+iSLEfHg8wPydlnGois5bVbIpD4ks1cqz9W5o6Lryhr9guKGRptxMUT2A8A8i/
SdZgfdGgxxDv6u1zEeajix+OQOmTWKWINTPPud0c3Lg=
`protect END_PROTECTED
