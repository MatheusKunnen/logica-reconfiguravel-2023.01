`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FTGDQpo+SXjKUmuOGfW52QheJ2wXrbXtUafUw4nz3qXt42TifAvbDF+0wBPvXwHh
1ybjHloGzrIwdh4nf0oTd2vSfAXGaOpr/0gWeqWQpIiuU4zcyvchBQZIlQ89UrWE
A14OdCsdWnkwK2Tz2RXahLufiWW7cqlaz4aZTRCn+zglOdSIhOV5vETbZ2IPwdz9
xiVGevilppGkemDx+QWNpz0suT1FN7UVYlJaDwCWUYbMFB7ffnlVhY6km5uZhr5M
IkwLMor74D/4I4+O9BDVJ9EIHuF70lmd3e8FpKvog/z5dl87sse/pqXvbACY5WFJ
G6KzNnRwerh68AGsWvKO7XyNLnmbAmZp/xi+lhQiEh8SE0ZgKdbcDEP4m0mMtLmM
I8FskHHxM/2nEwRiwuGdPKa8vifrC+odjIj535lQMhlWbRVxipnbdVwxLydNIxEZ
OgYh2votiU97RLv2A4dZXBV+RXsIJseDYo6m4f+5s09DSzLATRz/amS0LG5J0ftW
bXU2FWHmv6/jZyR/vSZ3XgchSci9JZ83Dmy9D11a+1QNHzZ0eCewcZnHQpWRa8mD
kPx5+tPzONN7VFEENFS6MGoYvoueCBHYzQNgxH0J37eCPpKHx+znpVhhh5/zmjz5
ON5aN83PolOqSlYOYYGNucJTwv2gzcTwtGNL2gZErGY1Hsg3MY7f+W0vPC2iyGaV
V4LJio2zxnlzgEyibPTAJ6TbcPo7NVrxi1zc0P63AqCkCAqV2v5/1/7ikw1ngMWG
VsUZaaaCRlAjDKQ1IaGlfcWo9HK5myMs9Pvtc1/4iqudkm9WjrdMVSn0aSPNB7YU
MN7PnAgk5sMAuQWBs39ot0n88Kjnp39V36fkMHInSKse6n27QDq+w/PU1UphAnAT
nKISrjQbT0TFB0KeRVrxG3ub/NnYG5BEkgcWz1h29aA1/4HS30KFN2qBpLmZ78uI
X2PF5M0LBzQuTWC9/bq7o+1zCEtUnd0b2o5kGA2mIVm2roxlM+V13vADTYtdLPtO
OD5NsSikxO7Kdj9WkpHrTze/JpYbOxK3Kni1H32tZZCOZI9wY/gBMaYw3GFZZXo1
0F1HEMa+8ahjXRtm4niY8tBshSgS8EyCf7zD8Vokt/WWZ3i54GNcPsEQz8mjVzNC
oJ6cuEtwJfN8CxMCDgHoh3SFTZUBefyQl8eZYJpkVh384eUTg5NaHT6SJoE1Osp+
hwiSG+LdK32BvKTEaPMGW3NSzKYaJsOxjFrPqGe0edyxC+nDiz1bWvXaAojXDvAS
iln+K5PxQIOFht9kV2ReEPy7Wd6J1T39OiX+R3QIrDuH9QTwtqdnyLusilQDI323
htMsENUiIZIkuI1B/vxuhZB18OzTP8b61iq75x7h+beJNBCuZe5RvwHcQdx0jIbT
ICms2qIF7p4wVnTuromDg007iMrsI/e7DHrXnbemXyKCmNguGt5DHuWWkqWaeW3f
qXLjIqj6WbeL+UsbZQ6xBnyKGgjDsOQ4btbfprc5WYjqtfg+xA3ctc4uXmmScO8Z
05YVTO5thg1yt4KvC6ZcbW1ddh1PAqm8BxFEfIX5r30zEePuibHdNvczlSF4JtSw
6ZwR8Qhz29aNhizIZKFTLjfpHrA8+5szYpahRjNDT4V4fIMCO9V5ywFDJTkiKd+5
Eg85PHcNuTLNzUW4S4WXH71a58TKY/VSX5VN0GYvhFVFxPVANlpTz3W9+UcM0tdV
He42YbszY7mTd6ArJtHLJKCsY0HhXk6eWOBGQnQHEJKfpFS7TDSXBiogLnUMiSAQ
FBg2TaDXM1xUvXlB1/BELOj1umWZjq7iWcH7elUTUGx4NrnxYq+pOVy86xG226a/
oFezyy0kNEnMT40V8dB3QqcdWN+LGERZIADKxkYyq/Q+mG4ZGrpVyZTijVRlxC4h
/uLnVMbjk2j+mbeUf9opzFZo5yFFkUwDeMrZNhfkU5fuP/b3+ZlZdVC9Rg3LrOym
ZDZAdz/JHyQ7eoc4fGsK8swudZnCelU5B1Ego/crhcl6GwFi/z8VAcxYGEhUYp+Y
`protect END_PROTECTED
