`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RAKCvlppNc9YlpOk3LWDd+AB4AkOHXilQa7YWIJ2NqH46/vGC2xza94qBDwkt15y
3GigdShpAVeYBv4uOqdRGXemidRiv/aVUOlxQygv4rjgMUpS+DWDZjgh0/Ttmeav
sMBcK0ICFP5IWo3NTvaCgLTNC09wtJUct51lWhV+t3qL2davnj+ToTi7ZFFiFBDn
2+eO2Rhv12TrG7EP+FBzM84mQ7rmrI5UWbQSTFL04GRKam8UnsjKo0TYS7OoGP/5
k6Aj5OHgFtBXS7QoheNvJF5SqMDIpRcQoIVhIIumfrRy06r7TBZPDIwOLeHthWSa
Jpz3fpiYcHfJP7illPpDE3P79u+B4YMuxigYPyJSy/9sU8Tct2bvo5hHyC7jj1jA
KX288VPayenv0tTmU6trfPRHzeZZ9Et+QaUJ0mdWZ2SNPjmKZjtVQWNXh5RXwBCj
tWNpvjLL7fv6RVqKmRme1bch2L/AREgzkO98pKWovHOel8C2V17uHADXH4UbOQ06
zQSQgtiCRKh+x3k+I3geVlC2Px+h8eCN9XKDUq+onbKwdcmQlBBwPm6Qc+IxA8VL
nAVwQlw/6cXLP7Zy6DBcvTayBLERPMJASBhIzK4rD38KPDgWgt8FPohqDcWYYZfp
g+F4IM8nhD8gpsWdpR1dLxdwSTOSQwPmS+durbIfeBOmdYmJ3NFGxYqtg4l+itm7
+WJieTit2/BBSGTnmPCvPPNmDpHqgeE0emGL3WfPuWPvlUFbOx1ZnXwYzmu1Jfbb
SvqSlhNX2Cd03qzcIP1ddiSk0Ukw8oeL02mM9OYGyQ0U0p941S/OBv7sepj9QyYr
bZLtzHMJHQZcQJDVT0YNFZuURqI/3o96VcQUXvsTc868ZqY4hGSKsrGar15hZi+1
8jkCeW2Oy6eJjFm+9pudOcNDv6B1Ubg1xPX2KPNn3FAz4eSbmSJzbR4z6HKKX0dq
eERnG5DuCt361QQn6ESqSRQ913Ngnw5dnnspDE6Xl8sID/Nq5aAUMldy8QPvqgjP
IMUe18ijhi+iuQtselWoGCJA0s/i1ldke1szm5E49Qtre25WnS4SWaKq90n9Q2ky
HtkN3Hh+ZeUW7lSCtmNttq8hUMGqxcnDnHVtzTwv9bxVjCn9FoMqxc6H0rSFsraQ
9aeiVXSWCf+ZKPGlknT4+xsAQJJWAyCa2WX/YMinl2IIhuEdVV76553hPF64wGq2
P2mvgw36G3c0T/CzKdEvj3zacTU7dD5FvsDjAgwk7WDe8jQ0cYf0VKBUpUyYoNoH
CKrKDSOdizk3D14f/vjveJRaO+lEPfI9Wa29av7TDy20faqwbm3st1jtkMhciocy
GCeMzbrqFsEAmAsz3zL6BCNSRhQ6pkodRZ3VWAXAOYNaUY1FyvkTY7jpq1hMYyfg
/5rz3VIwVB04Z/Bn1v9xq+u7Le5fE6TvD/gboJdJm5msyP+q95g5ss5Kf26WkIz0
JvfZz9GFKN9DwPCOY+w5be2VjCyXZ+F+tKl0aVAVI99fGZd1BsQXaIY9+3J0wjAi
3WzQe/zNlwu1Z5bhiG3ZIt4OEe1aMbDNABBZ0DqUqoiIXNXNRVSzF/FDzKXrj/Nm
1cERIZ2Z3VLJ7KCWOwqF4NIp+U19wHTBBykAdt9KfoapSWydTkhhNIMFNYcSic/l
BQBvSkRChtKMoaYdSSusMjFQ4TLNYl2Gh/Xped/v5NJ4gkxrx5777t88u0Ikw0P7
YqbdjjAC+rh3cXfLsNkFuyGOIWJQ7Fr10iOWU3ejM1crcxK6jY/djSNsfZUaFw2O
hgVWAVW9zaAENTslNwleTbOeKDmA5+hD6m6ILzby7LbHXmmFwJ3iwPkzpeTfYKoa
MXEUPDiGjvVVUREt0s+wnG3SHGa04JKOBfdgyHfveB184K7V2EDJ5xXJshEZOmyd
RaVJTduroQLxBi59Z5pbA+cwzEX5relSaUBRCzHV+/y3zTBbF6yKy3PGkAyjVKlK
UL13YmL687dpgFmL0hXpGEjrPnd+CTbtt0IInrv930gOmcRx+OvYCxkEu2RwGZg6
yiuFNqeUKJIFnq8nv9wxAxwfekgB4ZDjhzpVgRLGexNIctj0SglGSm2aob9t1dV7
vlL7G6sRPN3AoPSZzepSsE0GRcli1ra+2YUxp91KkxY+/h6N76w2q5nDtUIJCayM
b1KB3mhkcM7bfZyHDQHgZdFDDMRfVgH59CCDT/bGqVoeHX37jXaRKwvS8G4kfAWB
5PvesKIBkv3LAo5ZXx5Faw==
`protect END_PROTECTED
