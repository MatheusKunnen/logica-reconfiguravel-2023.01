`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ULkZOnrKF66+9GDuA0AeYDeMSYXXYXXhOEwEKMjdmC0Iz0S3/3P7uDDlJLEtMoH9
C1ExM2ziXNIN9KG3aKUzD03dwPy631Lx/H2eE6WwsHGbTsz8TzeghCBBywgkegSA
URo0/P0mracPgh2GBZtDZ1VdHVGoKZWaCoCxhbTg9ZI3JLReTeH/kxSb2rqwui9f
3yzaOuhTWydevvqfrAYPgC7YyGsnTw2qOcIWCzxgvEvveDx1dLM2aA1AvDn6g+KQ
xCqJb/E0VOkBcL4TeyNU3s9+tMciUN0LSjBFa6HdXHGMkujUaTLSXoK2mNDLfvlX
AqaTx4vOGI4VwA+iMIwFgmG2r7RjE5vUWhFHVYXbcKhllcOxWKI1wuq69rtnmSYR
z7QN+rbpvp7ctII/i93KBt0ccnW3mYvA50b6ep6Na4xZo0mcsqBfbxU242lCAkdW
JFVNHAy356Jlb4SGiSyUDycIo3Z9ZVGTWs/e86vxvbk7JTMRspAQHEs1H6Tlbr4x
J3NHNA/kIKf4Q5lx6vMRkg4XK1jMNkGeCQg7LRqaiuTdGUZa/rR4WO0bSab/q4Bf
EGcsBd6LDiW2uTGCAkzSgc0hr9Csm/S5oKZdAKpVxk4I5g+bLXLd0pMJEMJSYdIF
hmpI4K80T9dm5Pvw0ei3fMNv9IgORfCvaN0NQJTii43sY61rQ1FP8W403JcpBFQ6
xBtbX5W6mS9HHG9twKf4752VTN/aJSchwtAtNg7rawpEL98l7HZmjM4tEpzGO2bG
0v4RzjZCmHSiBMXHqi1da7UJvdMWBrh3sfT1DRQvfK9AWvX7y3+ajrTwb4oRlOdN
QybPpG+oNyKhlAd7tMvMa98QXllBt7ADArHgWkPj3UC5RAg9XxZpoo1MtVZMNBaX
Ltw3uob7RR7Lf756+x25XSLi/FvRhSRvP3f1U4Fh6ZRAGTP1EKm2D66RQgAH+ul7
qR8wXpS/udAc+9CqXc8193rC4k9frrz3xPv/Bn68uf2SLEtXyvLVVClXaAr+2gyH
KqRADj0ExkGv2tXT0quhe2b90sajx5qCsFBUbVszB08iqFUUf6ELrtdeTydPLl/9
5Y/Wp6udqdX6IRCy9RzkR+er/r05dNYrhdSEjsiPQPpS8vzzCqfpdc+J4jzV652f
KamgoI+eNC1W8FCLxkL4NzpxXvaA9JYJkPV1uuaeII7PQiCkqV6P+GDAI1aqcVBo
L4qZkKMgA5QHw8GgLIYDJ287FkDkAy/OvjRBup5+w0k9+F+s01zGS+2LW7ciR88d
8RuXsPTydXS+VHMBSvRwMqOLheFRj/37a5fmMv1462178khH7o+15oDgBtKpOpSj
Owv/RgseydzpsDQInW+LTdFZAsicMylgsXQC1vfvegQkGvdrtCxXDQd5R585HApf
5z/kbVmqfWW1sf4GfevOBGcftfEuswVWLQtxq6SPFAjWLJc2CSQSYV7PoMAZf2Au
dAnvGf9wuHkZfqLiOylR4h03FrybGis5/IdkDOLnHrGV818E5g1DJ/YB8lI5LjN4
PuWApo0U6I6UdQow15ZoZKJLyrndxrN/1tZdY5BcdQAr3KZQ9Z+Sl1a8i3DHz7Mw
cYrmdlb5hQAiN/zrGOnnJDkbDGOR/ueyuGkXs0S8WyB9GJGlHjdtFPSStltrk8Ub
35z0IkUKPG6MwpxfVN20TdjwYhDk4n1IFVTG4NzknnZCvX7GfKJboqaEyfm8p7ii
DtzVHI3mSYyonVSgv9SGRR+1a5Z5WAYsodHzxOrvSWshi2ugAwUFKIJhIuTmA9o1
O32PO8vq3pTnWDmF7TmoaUZnRfq5x8+K6J1ZT9reebF/XC0jpfFmo3zwWcEfU80I
F/gfiGmRbEMU6JfgPpY27DcWqzX6GNYU3sHQYKtibqQwHRXGrijrXaGwohnJkHKe
j9a9eR7yNidkLjKxIsA7+Psd8bb5fMwF6aN/F1gG5tdof6BqCxYGtQiMbdlliocN
N2j1PgzZLrtWdmBJvcd0/D7m2IlIIWB1JPtgmKjKRbFphlKeKMfwXCyqxOu0+xhT
`protect END_PROTECTED
