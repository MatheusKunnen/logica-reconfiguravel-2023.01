`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CWSdfSpMiVavNDScYdNVHCy72PJpa8BMYyblHu4TnnxBlT8LkVw5OKp/rZdAVJmy
3im91wQbfA2iWt3khdOQV7z4Z97LQpF1+5JzNhVwscJXDrEazPUPBR1iLfRCq99w
t/O9iNSoGiEQriyQA2IIVMNJWD8NpbNv2ZiQBKxuaG53qpVmTaSxa+OYzy7ZDTNJ
uHHcW5PmULCWvRbmNKDw+9JdjDJK/f2vInBLU7CSTRdwSQPu5YU1Wxpt0kC4LUUw
iVrEZ5/3nSiuw7gxYQJfggIdjK61gdaJqfiv/2Kism+bdaa0rz5ew+8Cp/hYSLW1
OXkK5rXx6QawbQ5brYNLbVR+JcHSKvV/fut/Z/LSwC4MYN0GF+rKO4xOUJ1YvJJn
GydxM45sAtpTGAa8V/TLZO44+iW2KrOPUjtvT9hqrc62sEMfWHU1jdWX1OPW0jWN
bc4+ansevc1ng6EITYVaPKHkUZ613HCgOful74QqxjxTUh1ks94o3x6k6yeKrIz7
sRiM/Rygw7g6r7NOfsm3kft+QoVClTNA8cEhqmI1Du0zRKmBitd0KplCjniBS+xr
AvOhUrYRsCUidz09F+SwAdXUEjsDAs/Iov11ZcCo6y7g8i2a930YA4FxOHeBfe09
HcIvPcZU8y92bp143fLIdHgMK2kZuEuXa4IpQV/CozTAHgUTazt3ZM2suigo2EvP
vwluCJOJZ9EUQ5EdwfAQTBvV9p1odAlkpSU/MEBCiDf+UxYwtUi+Poqh3K7BWgib
WchKoREEMd4piIeDbjxfstqiccxU/YWH+FCq3wiyZALsKzeB0s1Fww4yzAjCkBT1
EhywdhbAGG+/4ylgh0lkUbHUZHZspgW/UaCtUog4iYyxQTwRx2JPPEadGpNKbUwf
NaBrl4ZmxxWA5+Av/QQdhojVwc68zv+vBwmtMT2foGWc3KUlya/tl1910Si6+DI/
HllwxyZimFXNFM+aAFC/QgKIW7LZwQ+0GHOyW1wpw85gW9Spd56eoAqnhaQaLP/L
+I+Vi5i5wBEP0axdt0Bn44uJwNPC8Dl2uAfsR1AQThN1v6MOGuwVJEr6kwRNB0UM
xhtENEQuQy/vVH7uctKGGt8oAM1kvttCjUdJGrt+NtW6K+/q5vN8Tnmw4xn3ez+F
lMJj1mPlrVRjtVA2mDUb60+3SSFvFrwrL1Ni00NMzMz9++woORtoXef5NQsDJgw6
OKLtU/y9h0LZybSXrNosnxtSTaZV94vM3b9BvcUH5GaVB2huaXOpZ+wrb2yjL7OO
1G4HPrER7tW9gTko+MslQTwcfifsxaxjAhpqAc6iC6QtW/4N2gNOIb3X2JyygnNy
GJ95rKz3noN+Ixe2ikrVDblL0jrF8v24Pah0XT7Q3/dFw3S5MY8MZiC9KI/5j0lm
6gNtIKE7KV5sLwy7apEBXEWSZ3IImFsK3M0fxil2KV7Npim/51SA6mK5qDHbDHPp
odOJjKC4RHjLTibMoks1As7rCHLKK8TlmyKNV8ZDClcIExNTBG1m977qgTAtzf/Q
BzHHzud5LNPHM+/HZ0lKF9c2QWtWo9fN9GN36itDF9gnc83lrPoBgI3gXh8VspeP
7NyzfpyVySp0VrXD6NP3jM57X3DMzm3CweDIDerYjE6xkiHYbaEd0AnixtabAlyv
EOKbFSblbplcz9gBKngn2/uyESw2rC4w7+Omfji2Mku9lV3EJ+9pTkjrJejB/tda
DAyq/s58eCzjS8ac/AR6SKeYyE1sSHbD6BZ1W60K/PG2zSYaND3x7+Y60V8hS1JK
dhccO9nTcXQc7NEuwdcorMbC5E1RVWkj5fi5k78Dq4GuMEFhtOldiwNlGP2j9NgF
g7iYj/60EEytNkD29lH1Z864izaU3IA15+BH6NCPEapv3mzmom2vLUaQONkRM3iS
S0tpqiYw6lJ7b5zJRdH1qNT1eKnmF8w3sZXngjj8kHmJJXaWedyywdGcV8PQ441f
XoAXbWIybvIvvsGRuLJWw6EfWExHRjX4HAqJ4rudHDwm0yp7Eil5NHlhklCQo4Uq
T4dIV3HVUlWF2I6+Bb51NlBZGrkSbuXbxpjaTNvt2wc47+5W/JEs+HMzkyDnZvlz
xUpWtTY11t4RTt5oAQLPqTKKexgFy1ocxbijg0gKq+jm2WhzMt+nVI2uNUZyBrXw
sbZlgFye1kRRrClHz7g//GNZkG7zmSwwXqP4lfKyewu8m91FlKveOjfoDH1p11OI
emXY+/F/ucxZAM0tcGh4yurmTpeAw+aFswm9ZfjGYPVb9IXfymfz5iKqVTEdZuER
TV2r47Dyoeb+fWrR28kwlbiVjBempkuM8KYyBjum41GPNbHpXzNYsiqtCe1HSHCr
7CLA0Zn+pIlmIzwCdZ03FUWIYFNnL55yH0fSEkuu1FZfXoyQRNEvvnCkWm5ZrLRx
YCAlBVq+gkGf5PIQSXmiAfvXaHa7PEFvJqqSg2fbUzufZj/R4slQDIhrQ5jsBUp8
mKZD4LfWmeaUZWql4qs033oQqXD3/pBHIAIvuxQYxAlQcrnNb9jEz42aMkPAv++K
r1RStHbJieyyPCFQHVGe5+diOJglUjHo7dhcTsyl+fveXaboBQSUClTH1W6Gaaul
qSE8aYa/eAOzjMMq34RJ7FEsba+ampdpb3t2S/ieu19ESJEtPvmtxHkPhH2Dm21/
GdLxvOydY918DSqlP+n7VJ5GXO1hkaVrpEvvAK8ZUxtSAMKH7kwOcKBsY/5v01sb
v0LkryoqeALEE0kQAKegulyFgRPj6hHC2bJ1Ys4z7+N1xI04z9jslm983Px04GcM
jrpBZxCVvPEdOfarlHIhxUl59dzA7LUlRhwEEgsgSYV0vqfEzjKyOixJ494kQGN8
otOtw+Sbw/o6jeZMUjPsycY9t7ovZ3yiVhQFgf1SEEH1f+L3kSbGbRgvEwv09aCA
OLjvsFRfM2Senmz9yFXHRTe13ETLYTJEQdWbllDSPNedz5SJ6d0wXD1+m69IyASG
j+smthqmtaRckrJMIS2cseEdV3T0lq65w84MGKhesoEd6HBB/aaUSx1o1TFkbOpK
/LCO4ryLWmE3HIs8rnYhQQKUghDBJo6gZFpGU4cEt1iEku6PK4ZxcRZVg5xxC5ff
lo7HSv0C/OMR7cJgsB/oBjzN+qN1NMSLrOfF9j8z/u3W/20xAGrTmbLtK+HKqkqF
bAL33Wr6mvjb4EfLZKBFx/rH8Ok4UvBARx2ZbIS3GTy95ju2n7SipyAPE6pd43kk
/8aj2D3F2+Fs8lEaPmXbm/0ilSy36k9+m0wchFpHQ7PxXpeOPQhtGx5lBbHBBPr3
TDiq3c8fdWO6OvoChVg8TuOMHcYykaRlQE0LGhx+3E8Zu1M25U0H5swlXI0qbIRN
QodcKVc0kNXg51o9nB6zLAqVDqSRJ8yjd4gYTdhZVNiQd6/Ewtig+ODiZFd9O5U+
Ybhz6zGiZGT919ULb4BvG+VqrkH3Y63dRLUw3pUaJdZ7X18lm3LDFkW5aNG1+GKC
+ORQ0rtu80cdvOHlNhhDiUVEWautg61U84+9REJBurz6cNkcdA8YJKe0eatlLFwd
tRP7tKJMDSRL0hfTZ1jUNXGTZ4x6mzF4vHoBxDOQ8h/+NlAtsO7TafRApiC50GV3
LOSlrqfk4vE9NkdRQigX6xrqmTeS87prRzuxvvVD8ixG7tT/S5D2eN5SNokI6qXH
cRLj7cROO33StEeAENWF+AxxFzZE4O/LTi/wUXBorq4NYXWxo0BOYK1y9Ax3ALpo
6UA0eD2ih0arhpYURMwJrVNZQ5UJ3gMkAaJCTLm8YPG12ybJ1boUHWCRgd9+/LAa
IJgsbhNmVTEq96YTlYdr/ALQaoR6lm5P7mrwGrUW74QrFVEkphaN3tH6bPZdj5/C
brUu+V1uoT4iKlQl9rx6cV3Tyj+2jonDjyhEtAHfZ26EuXnD7B+llDcj/FeyH9gR
F7/EzNc+sWPmblGGSaJPPGoDP3Xklir70ylx4OQkc/vWfEao8cdFvnKnYjbmEMIZ
RslrdG+4fgI2XBW6EJzpwTbjXlq265baweoTsZEgh/XkI736ed/quHsPlZoe1Gu5
Zf6qSLNphcS5MEI2jMOpvWFG0W8gQnBw3dPHay2iGNuf+sgOJfI97s+RURh58LQ8
bdGHfgmbkHEmg5T9ArJIK/1yFTlmbgxsg+p9+8imF3MFnW4UCK4jABEFkpotDS5r
X53hE45kUN7IuBgLJyZZqSyzJIfwSfi3YKJQa99i3q7dBZzOu7wzkUxJwVp4+cZt
9l2m3oetd7i1wc3w5ut42jajzi8RRoAjt3GrlX2D3UN77C2xJk9Ua18KOPCMqeC+
ORa1BkBBUV68m8ehN/nn1KnZI9jl5DEx96D17gY1CgX3HGnfiCsWT5afDct7UTYu
P0CxgQHru2m3Tq58Z9UvlG+DxaJgwjY5OPySpa2Thfh8vXzIHktb83fgkxTqjrV8
5GTP8rZnYzW5TON+JNtQ5fo4wyRzUJBsXjqucjztyLYAIq94doOI6QEeCja2huP9
Hz5K3c2q5R+Muc5mDUW+vEqhXgkhRKG85lFresBEuhfbA/6YkMvw/NXWLgMftCWx
tYQVKpdKJ8IQqkTX/k0Sxvd41D3Z0zMK1qNDoNL2Hrk5M7ITlXhHsSHbm7B/N9yj
1TgsNLHW0jqpsSbTYXn/aCqg+ednPmu6fHe6mJuCxXUZPD4geJDCI+ZNRCGHM2hq
gXt1N0n2x7dBZif2W5f8C5Ov35AeY1rdkizPUhJXlWbHEDeo0D1vug9n7xomRtZu
c931gEKywvCVJ0f83wYqSq+C8+g9GUMj2e/LfwIee+bxeEOUhxuQzl3Jxh0C8SXL
0swU9Cldj+UlpSrIVCn0StIs1TI9TGV9g4twz3pHiauZDagGfpd4q2THQbWf/r8R
mpgjR21rg7ngrMzDRAJNjTpFaNiKiAjP5JXJ9ekpVb9a+4NRdaymporBgNKvIWI6
GW9kOySvQTcldyKS936HVxbZlFQ2lh8AFWyToAjt3kCtJfIJlzlw+c1eWZe1POIJ
Bc+eEK1AlZwvcHxli6G4BjOHgqZsOWkuwuG/mPU2RbNnntgSC7/4jd8nhVY2/hcZ
ZsvbZiwKmEacrFlpCcSNFkYkQ5Xa2YGwT1vlFFxhTrvMcPS20WDQ68Fq7a9Zjo4C
w9D3gqpC0xXjV8D3AdpXr9iZ0Vpqh8kod0aMorHjBfXv+6oXj+LO7o3TJ0nQDP2X
b9FFrTGeei9xINzhulUBHcEWzMPKjjuZgT3dmmOcUrTd4XaqrOqIOHI9vvSyu8Ue
vljBFIwkhPB4OZqlWlLXyc2ux6t/JQxZJrIKbuLlPtGPuWnLOyoMdbwJxBLTE1Js
YQGm1unfcJgo1u4oOEDrakGrc0hZSLCbjKgpxOo5YunrlV8e4Co0nQvN9cMjiyjg
uBSoPkSfYmTiIiCSa7OGmkPsECStrqqIbARPSqtY/paitsDxYpwW11v6fG6ir3b3
0LUGO/fEzRRnzJt9zfilraoI8fxfTbW42THc7r63wlgZ+Mb4wggKa5hZKTQS4Zgj
LkhXS+fuAMeTMKbzGgLgzsEfBCvq3nSYG4bfPOOKWiFyU94rqnvxEXiXay172vVG
yH9je7hA8s38bJhEfql8YrE+XPTOsJdMOVm2edwXgE9fjWYjqWDe8Yi0IxosUNqo
ZI70sjyamZmrqC2sjIOcc5Rg0+PFkkHUxei7aLrqq6to/4F1JzEhmPiwUjGMyWWo
ocsJMjikAKemJ5s1HqRnUoXbU3+YxwSRjFVZ3etzZqo5QQNlDz2ndrX2dVGfohQ5
vwzfX9wnGvyyoMCU4N87DQfIW+cCjGWVDreuaApgCqxPuin8tLKxTszMJiLE3z7g
UB/+b/v+kYsfbm5Px8uAXZkZMPaBEz3HSvABtx8abhgymIcSi+8dtv9BbDf/9MIs
a4XK4Go9bTwdupnkYM3AZGAsyvo/10nRBIVB0z3QdY7kvQfvuU+t88pEtvfph4l4
9tlyV/mQHOOfFlmmhcI3CLwRUN4Se7h9ruw+Zb5+2ps=
`protect END_PROTECTED
