`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ec3vzjzYYz0JxsnZfAErdDg3rFVRAClofmmNJp9d7N/fiOVjRu66A+T07TbyE96V
tz1JqwYhOSxgGI8DSHDU6T+/0lcdQVijpcEodCEaTsxQfhjaJrLIqoeDWtaasNYc
psNUkF5zHDPQABYdlpBOH/xwZcpcnZp4Tbs5oG37DMLM7WEDfThrYL8Wnf8i4Ukn
KqR+Uo27cln7FgwYeNhdJt1iIGhOaKPAxR1ejcum5puQGAzoT+sb33+67TLgM4ti
PkV2gnAfxxCLZShS5lBCzm7xpaGWIK8UiruUgDqXN7bJXI4dEcBf0UWyi3Duggv/
/fGM0wVdL6iAK3Yzgl6PiNS0uuyN9e3OIocCKJN9lZQ4klMw4lWIPQX76P22qa4z
2soD5at94LbzsYXHTmHnOjRNxhAfZODG1DW7kFtvVf+USHdFAjCC+nmhc1wc2hXw
QJeXihG3b1JUaDmrsjSZVSp/KFUTlxK1xRQYgvXO9sGoXrZr1zZ3uHsPXKieKtTC
XDYGRuilPN8dOj28yISYgu8i3MkLCiRaAnJt6xWNWmDujsn/9f4qQAXf1sRvm5dd
cfjkIkQp4nzwFOFrVuO7eArLC9h41JQRFceBXeHx3AEhk3tE8Cmyd380BAzPjoIV
7sNpV+8wWaxrY47ZOeAch1ou8TOwKkxqSvIx1IdLFr3PqZF2Mnpt5pPKhoX16CS+
l7adD44a1fMurI9Cmofz5ilF3e6s8X3cHs5th7GP1M1e2RYlFQ/HUMX+SqGUhEg0
MTL6Lg36vxUAekX+hjhs4oeNy6vNRr0CtLijlgkSqtv4x4/wTBTEyaDXCrG1bXjB
AlrlTugdJEvOWXfnUTlpV2vBSk61c4iRpu979WI9nfIvGwUqVoYVvAJ8WBKKFU5X
ruMcdDBwXuTxgvVmxE9R5XWgDuc0MR+kVjox34JUVZMVdzKaz4lBJXpjJjxGk/o1
uNPi/jcyoNZztUMoKTxOPwYkZoodk9tJNzMvAjHTslykGg56aS5b0Z/Rdwp5TRu4
/RZY65EUD4u7QccAcYV5AvszS/5Z2N7B4HCAk5UNb9TbOE2TuMzOH+Qt+RWTfS+E
0HyQG1f3+wNt6sfQ9UMIpPWaBUHoMR3SS0npR0uJL29/RPsN0uH2ZaSWBCZwV0V+
J6gVhgFqCwHTFDcT3NheJDM+pNYhjbue+KPw6DWg1glBOubmi2ZslXd/4G2Q3Teu
RUnfbNSwYmfUrxPt8iFYepIhRmXVOOzmMb0IEtBtxIYRznlmp6ky1LFFNqEcD5P8
LHvwt51+QNNAazoe0cvYiueQnvvDA4PajahLW8molUAR+/3+byY+8pjPW2+w751X
1f+7QikZk60CgQUw5yhusMN59N3aLHDGgKsXpQtr5Ey9ACEhpH0iOdiC5qokaZyn
9DsysSw6hJHdXSCkh/ySw7kVAbOza3tFE4GW54wpDV3i0MNBxXgAFVUrv0kzLOp6
+lEcAvmJsINObdn/Smjgx97pf2zFkzcH/4jeuMS+pMFlBPtlh2nMOBVrWdxgd+At
Xr15qhpuksjiI32f7OidUhbxWopHregrdOcpH96NZR8GEnaMXOey1zaKm44i3ORJ
e6zxmQ3PXVYAfohzm/xdrxQMxvjnuII/w3pOpEwV5ZPIj7i2FgeZZvhtj4J3OAG3
lWh0KlFoNJofZL6PeNEjMZqFPMFbTgPVC6XrjTDKEVQpXGBohuxGPoWDOM8UG5bt
Gi29eqLedQ/1hWRORmcPlSJE5ZrV+acFd08YixWbWb8vX1V3tV04/DLOaC+7Qz8D
tjN9Mc6VWlZ10A1DGSXsh9BydVDOpSbsWs04Ltb7LeUyi/tAQLsLRDVJaO8MrgBb
um7FvyJDynzLsKX8Mw09DJpMk32tzAUsOD1oA7De40A1YRlnk/Ed9O+XmzuXApVL
sSMNeCwT6NCGgmN2UKdGo0jVsNunHwRjEr0+ppl9o7fsErwdon2qdzNx+xYD2mx0
WbTvw7yq+3lPplf/sQ67Hg==
`protect END_PROTECTED
