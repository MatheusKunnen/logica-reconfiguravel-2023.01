`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3KjpGaQctbpAmpn0oRG82De0GYRWB73Lmab7L50WRVGaZVxhp9G2CujdsLNwIhJ
T2cw7VpzQeAOhSMyVpw1sL5KONhFEBlvwDbLMq7u7DJBhVuOjilcYqDh3J800eYw
bgD0+5g+f8kxAVLML7soh8xUYQ/P0ERmztHX3VOWyxm0v0Zmkix4Xe+GAp/Spl05
PmyitBUtkcjWFC8XRxZru+kWmKqlI8/R4kYxnCpvo6A9P0IMi9CsJLlwcEujLcYO
surSiUYml3ibjhTEMC4K4SLiaHgmWgjLcAFpO5nuLyFyWgQz1tUR/l6aRyZ/7mC7
sMD6BjjCnrZiPXx8f/2vsnrLD2607i26aVhevCFo4KKyrBm0qAgYXFcFMssmHN2+
QCR7ekzwFed7lPO880WL64552Cb1HuevCbwsy++YG4JQKZzTL2ekXwWb5GL3PTSS
Xrs1w+8MtdQdzkvg+fRdDqmjvVNWrDA1YhGHc63dKtd4Zu1i9Hordj+hENDVNDLr
BLx2RCIWm3yvcYdUvByP2DnZIhWCHZN5dT9BOpl/uL5vR+1+hGvGXFzYOe7sBhLo
X3tIlxKueKoPx1pZ7C0ogso/hk+vbTY3o4EBzxaUpyLIiDejkMTLugGWvUDADbcG
dGqDGP/w7Kr4OqFa6Kjhzi1uSg60OhMgVbjnsSr7gw/VpHhcyow+cklH0iATIBR5
EyIeCV5Q6tRqVLx1iDEeL1Fy7484znIogUgd8wsnyM3lN6jVaIotWA1EtUMfve8H
qAk1JQYer12QsM9mpQvc1jKC9iLIQhR64dm48kfSs7M6RVrDkxnUiwF0s3DIgYpk
zsVGjVG0uujCZhhOVrGPUf9SY47ChZWgIEKviUegWE2srxpcOSbl0y5MHccPGVvI
8JeNds9+jCZwMoTSUmmC13JscmhiEuKKlRfZf/HTB93blgqMKe+W+nNI1snP09F0
bNYh5wsXKML4Xo4uUF9dLy2VivKKITeRXL0vuvV3VT/A5lKvnu5c4+3AJuyw/vkX
2XTLKFqYzOw3h+71QdsXp/5XQ6meXpWA7vUSH4q9zgUcR/Bp/UUq5nXk8UlmywNq
dFp6GHFkfM9S8dumCoZbm5Uolw8prgmduqDmD7acLJpsp4+axdchnNQmBfL+dGd0
WCOPSXeeaEGO7eLnQ8nCyqI0QojMsqoMT6PKJ8FPiGEWGo6pzRBSXbIzN1FOltm1
lY7LEBDUbYgZJtPLxFEBlv7VWUWei9/Ugp9MrKxqFCNkL0aMDyOcEdkn6qsHh/I8
EBm/rsIRy3nd0bwJleVqIniveUcJz3YcJCQLBtX1BTfaP2DHMZqotawcAVEOMlS9
soqUVVre9ocnJS1l5kkECA8IFHPKNWN06vIShVBgAAUs2IMz8rPesJGv0x4f1UxQ
v4RZUIxtjIfvuJvbX+z1Yv7ya0WNvlsx0ZsojpErkQJY0r3Itq3U5dX70E1fXM/b
dEzuc1kJkh5qdrC6n/vA/gQtLhBGZ5qsSis5rEixbh0FEAkjO0w6y612NGlNekRX
cyZI+9d39lADjRm182sb/84yGUcYyKM6jv/2UTpMDESSSk1VPNQZs3xNA8hHoKDC
L8e5zGQSDaZPAtcEb8wUWQDmU4Y4ifv+izRTg29Jz1N0/SqdaKVvt8ljpbr2eftW
opKrorXiA8LhhUbqUXUSYBqDrM5HfAPdJdqjlgGsc154Hp2Kj2vvgwuPOmXz18Li
LRKq/kTlUDRgtuBEvIIJvS62kSdjZERZJxixRa+NrzhI7faZdtMHxP+kyWXxE+Zk
MdUUO8x7vxWFCpcoLFcWidnDAcZQnshAK3gRzgb7zyH42KjpuefC8EMLaIrOICsi
KV5SpXVTUikqqcX5oxMjeabICGZ1opd7JlywyFD2d2j8v+CMlgbMlBBMt88CVchD
QMzNRLcq+bqSghwXe5wuGRmgNfFy83Xl8HdsItfAVsF4fjjTECRQXyGBH3tc+aRu
wqaYJZbGPXkG06qWWune1z/BBCi6Vxc6evpBLhg3ZjGpeF46w8bXhdGw8Z52AybE
AXehqeHcsus7R2f2nwlJ6529mCODHN8J0TzrryVPDQ37Q7cKNtbE53SZ6CrKuLzb
DIyIuWwB+PFCpSv3ispAYAyy1Lx8wKxPE3/mFwiKLWthoZE4pFrZ3orF1NL656Lb
4+a1ZqSjaMSEtKBDmTyCKyoaqPC1X1qQ5ptwHtovpoM5lYBjX1FJ4PGx9nGAChB5
rcaX3tDDrLAZW2/kiHjaj1Obj5qF7AwwpzvUrEAeCcFy1ILEVQ0nsuSTEZeH4IAs
DzWFgl0vefnoEFO5vEVIKimkKKxiFrguFC9J+7yhZN+Gpod+j2CgwgfSHrKsxmN5
CuYi+OI/lz1H4R/FqiLudjc2hiKAw1tEGUmmWFEuqpph+MbsC/Fnxrt3Nlvyn4gC
OoGAzKCpOc21qT2z9dJrSxkj3e4Rr3R+F2S9Q/jQqUVJ4ewaHUo0l61kbNufra5Q
aJsFtmJadgnz1PikhwhBcUBxRuN3Bdytrrw3ycsqdtyZnLzwBz7qzyfHOYvb7H1i
7JSI9C3Od88QzgbGh4/AjFZlBhiZhuykycatePDWRafTGZc/b68KfiGEUEo2r9K5
4PiHlqfcwna9OqW+beo9Mj7hKIdZzFcoH/Q3KauFNBb1BeB6vfbpVySJLTzYNltD
dUi8GJpclC7tGXCqOV7eYPpMUQzCx/XeWRsHOxYx1sQQNQohv9RlrWHUXz//dmu9
AnAADVJLcBIQ0D3o9+wK+otwMYHItG3Iyvx4CNG3mj49VvUiSkaVUplDSInxOcOa
PNzdQpI3OmiFXAyCGNc7WbvHyCXqT1eunurqxuPEdD0EihPLOYvTRP4HEG3Bjr9y
V7mxJqUAg6dchnLFR0Jp95f2XgLqqDt0fKivooztmm9pbwIgjr1QxK2AuKwZNWMD
e5EkCj42ArB7KyFVT9tk29ODPqTYr4oeEMM2Ql3uAWRTxtN1t0Un+jLNcN1de57Y
JAqdK4vNcDHtKA2xe5mow4IiGjOBklQzUN0udsSoQhzT+nY9Mq4yfI89mKmjChVt
8/i7wRjb4hNidmkgg89Yjd9HASwamegCZGhoSbTtd0HhOrooyYTXi3Q95YjNo+VZ
cjZ8acPlzZpYcqI5TBhTFmWtsTofI9/xHQK/L98wMH54Bp2XYUbH3r10+wS0LJvS
Z21kHKDuWtV5RLYQpbE9IFB7mCOuTHq6FQzwvvOrUdyU79++/se9ciRgpgfKIbeP
aQZ2diAFD7ZisD3YsJCN1BrkoRV1F+gA1a0Dv2ixB3m4qxFnvKzRik40v5INdkkZ
TiqZVB0t/SlLScGLnn0bxyb6YRbVtxsz7CC5iqHA89aV+IBnIhZO9LLRrh2Hbp/f
fomnmz1mUx7mHFBVt1x3DAQMRmuDR3YTGzVMIHl2eua7yD7e74YNr1mSWP+U4Cdc
gMdBuGDtpfrW1wb+LHByK8rFPsyoYZtBkgtQ3IeRWvuD16TYGWTMvrTVu+bgihBP
ePPDxrnR8YUe/95gyxUzHzW6mGB6FIy1uVVGB6fOC7P2G29Eg5l/9XB6ZZZSbcXn
W3VFkMrq++690i6+SwDBxQnR7cEKPhza8L1QGmwdsgjgPtHxYxToFL3CIQ0cgq6t
0SlrfrAVeBRVgKJr/U65Kk9N2nudEMusrz+q9v0qlYeJXB6oi+oY6BpvmJhOWBN9
bsvDDHFnMcGRUg4ct1sSdVMvCY17J21tWEBvc0LypVzA1XX9iv/hLf6oCv1ww7R+
gF7D9GRWEmSC2t4nz54Wp5YwoxhAedfwtQM+HwbyMN9z+3GZaR52fAIkzB4fdOVp
IS2z9m9s4NvkN57Lr14QTN90eUjJ42LEtpOC9UumC4RmPpQRBNH6yuqxey66B0xv
J7Jv0v1pDCOjqk/PLyKGEgcqchaeaPCpHpYFUsPUG8h/lt2hYGv2U/2sdZKXvliI
1crZAlRK3M/IkaXT523XPPuxB+nMn35aF+9i206ESIG1CEeZrMpCSQ03t99Je/hQ
6RnOnCwALt0DmuBtXTujgw8eYPLZjGcQ3KUuaOTcnC3NCRg0fdKUQI4yMmClLhwp
sOPQq+yhGvc5/ewtQTkpjux4wyS+ygOhlMy7CJPc3cyexCgrm2oxvinsFnjg+ONo
30yKcWs2VwQFowXVCVWzFiYFe8uKr6APWAk36W1Y2UmSKFL4yEoPp2asUNboduCh
mBfyNwEPXTErshZLc3DrpKawrEqytfVBSJ/Q6DMGdykpc4GJDTg4/E8vCKVklH0W
LcfTOGx1kxITajpQ/UmBinoq1gr0NwPb4tv6fumts0XC4Uo5vfKlOf/E3Tlluzd1
BGu7pitfV9BQzkbRL99k8Oglu1B80GMb+uMeucgAKPp3gVsRjNyd4BkIL334bNhw
aOr+Mv2FtdzVZ4U4JSs1OOAPdhCtRn2viFmOb3ojZTmkUuwmNXX9pS9n9dqJaens
1KExMKVNF0kesFT02IwhbVvlcK+2svILwthkiiQv0M08DvUllxaO4ActKuYXCJKd
UcQUbhquHjO3WTouaET9voLsi58MUPXPjOuhhmb0MwLbZPKMHNAQSR5dSTkEbMls
SfPKfH/E5wET4OwIuPYmAcxc2mJ/7BQmmtC4WFowGgy+g78kqLtLnI2Z4NPOS/q4
p8rk8kw3y5pcwtehq24a9WmK7qsJtmSF8yqEXNKhPYxcJpVpXOGJ3T+QB2m4/3hP
14vm/pikKJ1A+hoc/IBWLgFtFpP1BcTBhU4mxiqCweU5CVOMC+D8zGY+uOFCHMTN
VvAAeDjwSndwYZeZuM2ZBF79BuWNYRJoWRlR89HqBAvKc4yAUU39Dgp7KeS7srfy
4O4cZuGYtOAkHxbRMgYE6xCwe2QMrdFJP2Qs+B/9phOcy8NRjWVoNUQjYlszXlTD
O+HnxRyW43gPGf2a+UcBeJpv5wOiuBudajLkmErMUgx0haTOeOhIvHlqwGb9yyt0
vMfKYgMbo4fBCzjRKo5mEamssXqY+7pz0t4lFjPl8J6P+EuIcPhZV3QjNu9xY/s7
hcvXOHz212R/EPeO10Hc1kLjZTRIWis0Klpr6KCiJ9izn4vtg2UrijbGBd99hTQO
vmCG9h30X0U1qpIPJNnXiqM377XSDOT+vyvmwqvtaxeIKdSNSxqulJBs03OI7GLr
qf69FlclS9M1/y2hUod68HVAgfF1ed4+xSXhPOx2e1Rvd8omHLTnkMy2vGmGrut9
/GSOXFQTyWkcFOAwgrkZ8iUh3UpJMWn5POwMMCgdlx8ow5mZKjeBA8op++AkggHg
cI2ygaO6zYb7+3nwPaROrJCrFeuAM/K7PJgvcgtn3iO2h9GrrgLOULvX2eMoDC7/
6wnjs29kUAlHZ65KVp5y2JFw3oWQSuQ5CxrnqiIA6Z/0D4tr6gPBPw2kH6ll5zoz
CqJ7vXex/eqgV31ene92z5h2Y5htdUIhUGSXgXzbjqz6mzSikoQalVvcVWZP5Mdi
rW4LF/VZNW36n6iIXeTBZg==
`protect END_PROTECTED
