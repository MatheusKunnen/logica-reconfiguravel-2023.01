Library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

Entity BRAM_tb is
end entity;

Architecture X of BRAM_tb is

component BRAM is
   PORT(RST       : in  std_logic;        
        CLK       : in  std_logic;        
        READDATA  : out std_logic_vector(7 downto 0);
        WRITEDATA : in  std_logic_vector(7 downto 0);
        WR_EN     : in std_logic;           
        RD_EN     : in std_logic;            
        CS        : in std_logic;           
        ADD       : in std_logic_vector (9 downto 0)
		  );
end component;
signal GND, VCC: std_logic; 
signal rst, clk: std_logic;
signal READDATA, WRITEDATA : std_logic_vector(7 downto 0);
signal ADD : std_logic_vector(9 downto 0);
TYPE state_type is (idle_st0,idle_st1, write_st0, write_st1, read_st0, read_st1);
signal state : state_type; 
signal INTERVAL_0, INTERVAL_1, counter: integer;
signal address: integer := 0;
signal CS, WR_EN, RD_EN    : std_logic; 

type mem is array (0 to 417) of std_logic_vector(7 downto 0);
constant data_nomes: mem := (0 => "01010000", -- P
1 => "01000001", -- A
2 => "01010100", -- T
3 => "01010010", -- R
4 => "01001001", -- I
5 => "01000011", -- C
6 => "01001001", -- I
7 => "01000001", -- A
8 => "00100000", --
9 => "01000001", -- A
10 => "01000010", -- B
11 => "01000101", -- E
12 => "00100000", --
13 => "01010100", -- T
14 => "01010101", -- U
15 => "01010010", -- R
16 => "01000001", -- A
17 => "01010100", -- T
18 => "01001111", -- O
19 => "00100000", --
20 => "00101011", -- +
21 => "00101011", -- +
22 => "00101011", -- +
23 => "00101101", -- -
24 => "00101101", -- -
25 => "00101011", -- +
26 => "00101011", -- +
27 => "00101011", -- +
28 => "00100000", --
29 => "01000001", -- A
30 => "01001110", -- N
31 => "01000100", -- D
32 => "01000101", -- E
33 => "01010010", -- R
34 => "01010011", -- S
35 => "01001111", -- O
36 => "01001110", -- N
37 => "00100000", --
38 => "01000001", -- A
39 => "01001110", -- N
40 => "01010100", -- T
41 => "01001111", -- O
42 => "01001110", -- N
43 => "01001001", -- I
44 => "01001111", -- O
45 => "00100000", --
46 => "01000011", -- C
47 => "01000001", -- A
48 => "01001101", -- M
49 => "01010000", -- P
50 => "01000001", -- A
51 => "01001110", -- N
52 => "01001000", -- H
53 => "01000001", -- A
54 => "00100000", --
55 => "00101011", -- +
56 => "00101011", -- +
57 => "00101011", -- +
58 => "00101101", -- -
59 => "00101101", -- -
60 => "00101011", -- +
61 => "00101011", -- +
62 => "00101011", -- +
63 => "00100000", --
64 => "01000111", -- G
65 => "01010101", -- U
66 => "01010011", -- S
67 => "01010100", -- T
68 => "01000001", -- A
69 => "01010110", -- V
70 => "01001111", -- O
71 => "00100000", --
72 => "01000110", -- F
73 => "01000101", -- E
74 => "01001100", -- L
75 => "01001001", -- I
76 => "01010000", -- P
77 => "01000101", -- E
78 => "00100000", --
79 => "01000111", -- G
80 => "01001111", -- O
81 => "01001100", -- L
82 => "01010100", -- T
83 => "01011010", -- Z
84 => "00100000", --
85 => "00101011", -- +
86 => "00101011", -- +
87 => "00101011", -- +
88 => "00101101", -- -
89 => "00101101", -- -
90 => "00101011", -- +
91 => "00101011", -- +
92 => "00101011", -- +
93 => "00100000", --
94 => "01001100", -- L
95 => "01010101", -- U
96 => "01001001", -- I
97 => "01011010", -- Z
98 => "00100000", --
99 => "01000110", -- F
100 => "01000101", -- E
101 => "01010010", -- R
102 => "01001110", -- N
103 => "01000001", -- A
104 => "01001110", -- N
105 => "01000100", -- D
106 => "01001111", -- O
107 => "00100000", --
108 => "01000011", -- C
109 => "01001111", -- O
110 => "01010000", -- P
111 => "01000101", -- E
112 => "01010100", -- T
113 => "01010100", -- T
114 => "01001001", -- I
115 => "00100000", --
116 => "00101011", -- +
117 => "00101011", -- +
118 => "00101011", -- +
119 => "00101101", -- -
120 => "00101101", -- -
121 => "00101011", -- +
122 => "00101011", -- +
123 => "00101011", -- +
124 => "00100000", --
125 => "01001010", -- J
126 => "01001111", -- O
127 => "01000001", -- A
128 => "01001111", -- O
129 => "00100000", --
130 => "01000111", -- G
131 => "01010101", -- U
132 => "01001001", -- I
133 => "01001100", -- L
134 => "01001000", -- H
135 => "01000101", -- E
136 => "01010010", -- R
137 => "01001101", -- M
138 => "01000101", -- E
139 => "00100000", --
140 => "01001101", -- M
141 => "01000001", -- A
142 => "01010010", -- R
143 => "01010100", -- T
144 => "01001001", -- I
145 => "01001110", -- N
146 => "01010011", -- S
147 => "00100000", --
148 => "01010011", -- S
149 => "01001001", -- I
150 => "01001100", -- L
151 => "01010110", -- V
152 => "01000001", -- A
153 => "00100000", --
154 => "00101011", -- +
155 => "00101011", -- +
156 => "00101011", -- +
157 => "00101101", -- -
158 => "00101101", -- -
159 => "00101011", -- +
160 => "00101011", -- +
161 => "00101011", -- +
162 => "00100000", --
163 => "01000111", -- G
164 => "01000001", -- A
165 => "01000010", -- B
166 => "01010010", -- R
167 => "01001001", -- I
168 => "01000101", -- E
169 => "01001100", -- L
170 => "00100000", --
171 => "01001000", -- H
172 => "01000101", -- E
173 => "01001110", -- N
174 => "01010010", -- R
175 => "01001001", -- I
176 => "01010001", -- Q
177 => "01010101", -- U
178 => "01000101", -- E
179 => "00100000", --
180 => "01001100", -- L
181 => "01001001", -- I
182 => "01001110", -- N
183 => "01001011", -- K
184 => "01000101", -- E
185 => "00100000", --
186 => "00101011", -- +
187 => "00101011", -- +
188 => "00101011", -- +
189 => "00101101", -- -
190 => "00101101", -- -
191 => "00101011", -- +
192 => "00101011", -- +
193 => "00101011", -- +
194 => "00100000", --
195 => "01001010", -- J
196 => "01001000", -- H
197 => "01001111", -- O
198 => "01001110", -- N
199 => "01001110", -- N
200 => "01011001", -- Y
201 => "00100000", --
202 => "01001011", -- K
203 => "01010010", -- R
204 => "01001001", -- I
205 => "01010011", -- S
206 => "01010100", -- T
207 => "01011001", -- Y
208 => "01000001", -- A
209 => "01001110", -- N
210 => "00100000", --
211 => "01010110", -- V
212 => "01000001", -- A
213 => "01011010", -- Z
214 => "00100000", --
215 => "01010100", -- T
216 => "01001111", -- O
217 => "01010011", -- S
218 => "01010100", -- T
219 => "01000101", -- E
220 => "01010011", -- S
221 => "00100000", --
222 => "01000100", -- D
223 => "01000101", -- E
224 => "00100000", --
225 => "01000001", -- A
226 => "01010011", -- S
227 => "01010011", -- S
228 => "01001001", -- I
229 => "01010011", -- S
230 => "00100000", --
231 => "00101011", -- +
232 => "00101011", -- +
233 => "00101011", -- +
234 => "00101101", -- -
235 => "00101101", -- -
236 => "00101011", -- +
237 => "00101011", -- +
238 => "00101011", -- +
239 => "00100000", --
240 => "01001101", -- M
241 => "01000001", -- A
242 => "01010100", -- T
243 => "01001000", -- H
244 => "01000101", -- E
245 => "01010101", -- U
246 => "01010011", -- S
247 => "00100000", --
248 => "01001011", -- K
249 => "01010101", -- U
250 => "01001110", -- N
251 => "01001110", -- N
252 => "01000101", -- E
253 => "01001110", -- N
254 => "00100000", --
255 => "01001100", -- L
256 => "01000101", -- E
257 => "01000100", -- D
258 => "01000101", -- E
259 => "01010011", -- S
260 => "01001101", -- M
261 => "01000001", -- A
262 => "00100000", --
263 => "00101011", -- +
264 => "00101011", -- +
265 => "00101011", -- +
266 => "00101101", -- -
267 => "00101101", -- -
268 => "00101011", -- +
269 => "00101011", -- +
270 => "00101011", -- +
271 => "00100000", --
272 => "01001100", -- L
273 => "01000101", -- E
274 => "01001111", -- O
275 => "01001110", -- N
276 => "01000001", -- A
277 => "01010010", -- R
278 => "01000100", -- D
279 => "01001111", -- O
280 => "00100000", --
281 => "01001101", -- M
282 => "01010101", -- U
283 => "01010010", -- R
284 => "01000001", -- A
285 => "01010010", -- R
286 => "01001111", -- O
287 => "01010100", -- T
288 => "01001111", -- O
289 => "00100000", --
290 => "01000100", -- D
291 => "01000101", -- E
292 => "00100000", --
293 => "01000110", -- F
294 => "01010010", -- R
295 => "01000001", -- A
296 => "01001110", -- N
297 => "01000011", -- C
298 => "01000001", -- A
299 => "00100000", --
300 => "01010010", -- R
301 => "01000101", -- E
302 => "01001001", -- I
303 => "01010011", -- S
304 => "00100000", --
305 => "00101011", -- +
306 => "00101011", -- +
307 => "00101011", -- +
308 => "00101101", -- -
309 => "00101101", -- -
310 => "00101011", -- +
311 => "00101011", -- +
312 => "00101011", -- +
313 => "00100000", --
314 => "01001100", -- L
315 => "01010101", -- U
316 => "01000011", -- C
317 => "01000001", -- A
318 => "01010011", -- S
319 => "00100000", --
320 => "01010011", -- S
321 => "01000001", -- A
322 => "01001110", -- N
323 => "01010100", -- T
324 => "01000001", -- A
325 => "01001110", -- N
326 => "01000001", -- A
327 => "00100000", --
328 => "01010010", -- R
329 => "01000001", -- A
330 => "01001101", -- M
331 => "01001111", -- O
332 => "01010011", -- S
333 => "00100000", --
334 => "01000101", -- E
335 => "00100000", --
336 => "01010011", -- S
337 => "01001001", -- I
338 => "01001100", -- L
339 => "01010110", -- V
340 => "01000001", -- A
341 => "00100000", --
342 => "00101011", -- +
343 => "00101011", -- +
344 => "00101011", -- +
345 => "00101101", -- -
346 => "00101101", -- -
347 => "00101011", -- +
348 => "00101011", -- +
349 => "00101011", -- +
350 => "00100000", --
351 => "01000111", -- G
352 => "01000001", -- A
353 => "01000010", -- B
354 => "01010010", -- R
355 => "01001001", -- I
356 => "01000101", -- E
357 => "01001100", -- L
358 => "00100000", --
359 => "01010100", -- T
360 => "01000101", -- E
361 => "01001111", -- O
362 => "01000100", -- D
363 => "01001111", -- O
364 => "01010010", -- R
365 => "01001111", -- O
366 => "00100000", --
367 => "01000011", -- C
368 => "01001111", -- O
369 => "01000010", -- B
370 => "01001100", -- L
371 => "01001001", -- I
372 => "01001110", -- N
373 => "01010011", -- S
374 => "01001011", -- K
375 => "01001001", -- I
376 => "00100000", --
377 => "01001000", -- H
378 => "01010010", -- R
379 => "01011001", -- Y
380 => "01010011", -- S
381 => "01000001", -- A
382 => "01011001", -- Y
383 => "00100000", --
384 => "00101011", -- +
385 => "00101011", -- +
386 => "00101011", -- +
387 => "00101101", -- -
388 => "00101101", -- -
389 => "00101011", -- +
390 => "00101011", -- +
391 => "00101011", -- +
392 => "00100000", --
393 => "01001010", -- J
394 => "01001111", -- O
395 => "01000001", -- A
396 => "01001111", -- O
397 => "00100000", --
398 => "01010110", -- V
399 => "01001001", -- I
400 => "01010100", -- T
401 => "01001111", -- O
402 => "01010010", -- R
403 => "00100000", --
404 => "01000100", -- D
405 => "01001111", -- O
406 => "01010100", -- T
407 => "01010100", -- T
408 => "01001111", -- O
409 => "00100000", --
410 => "01010010", -- R
411 => "01001001", -- I
412 => "01010011", -- S
413 => "01010011", -- S
414 => "01000001", -- A
415 => "01010010", -- R
416 => "01000100", -- D
417 => "01001001"  -- I
);

begin  

INTERVAL_0 <= 10;
INTERVAL_1 <= 15;

GND <= '0';
VCC <= '1';

gera_rst:process 
begin 
	rst <= '1';
	wait for 15 ns;
	rst <= '0';
	wait;
end process;

gera_clk:process 
begin 
	clk <= '0';
	wait for 10 ns;
	clk <= '1';
	wait for 10 ns;
end process;



DUT:BRAM
    port map
	   (RST       => rst      ,
  	    CLK       => clk      ,
        READDATA  => READDATA , 
        WRITEDATA => WRITEDATA, 
        WR_EN     => WR_EN    , 
        RD_EN     => RD_EN    , 
        CS        => CS       , 
        ADD       => ADD       
		  );

gera_data_we_rd_add_cs : process (RST, CLK)
begin
	If RST = '1' then
--	   READDATA   <= (others => '0');
--	   WRITEDATA  <= (others => '0');
--	   WR_EN      <= '0';
--	   RD_EN      <= '0'; 
--	   CS         <= '0';
--	   ADD        <= (others => '0');
       counter    <= 0;		
	   state      <= idle_st0;
	Elsif CLK' event and CLK = '1' then
		counter <= counter + 1;
		case state is
			when idle_st0 => 
				if counter = INTERVAL_0 then 
					state <= write_st0;
					counter <= 0;
               address <= 0;
				end if;	
			when write_st0 => 
				state <= write_st1;
				counter <= 0;
			when write_st1 => 
            if address = 417 then
               state <= idle_st1;
               counter <= 0;
               address <= 0;
            else
               state <= write_st0;
               address <= address + 1;
            end if;
			when idle_st1 => 
				if counter = INTERVAL_1 then 
					state <= read_st0;
					counter <= 0;
				end if;	
			when read_st0 => 
				state <= read_st1;
				counter <= 0;
			when read_st1 => 
				--if counter = INTERVAL_1 then 
					state <= read_st0;
					counter <= 0;
				--end if;	
				address  <= address + 1;
        end case;    	
	end if;

End process;

process(state)
begin
		case state is
			when idle_st0 => 
--				READDATA   <= (others => '0');
				WRITEDATA  <= data_nomes(address);
				WR_EN      <= '0';
				RD_EN      <= '0'; 
				CS         <= '0';
				ADD        <= (others => '0');
			when write_st0 => 
				WRITEDATA  <= data_nomes(address);
				WR_EN      <= '1';
				RD_EN      <= '0'; 
				CS         <= '1';
				ADD        <= std_logic_vector(to_unsigned(address, ADD'length));
			when write_st1 => 
				WRITEDATA  <= data_nomes(address);
				WR_EN      <= '0';
				RD_EN      <= '0'; 
				CS         <= '0';
				ADD        <= std_logic_vector(to_unsigned(address, ADD'length));
			when idle_st1 => 
				WRITEDATA  <= (others => '0');
				WR_EN      <= '0';
				RD_EN      <= '0'; 
				CS         <= '0';
				ADD        <= (others => '0');
			when read_st0 => 
				WRITEDATA  <= x"00";
				WR_EN      <= '0';
				RD_EN      <= '1'; 
				CS         <= '1';
				ADD        <= std_logic_vector(to_unsigned(address, ADD'length));
			when read_st1 => 
				WRITEDATA  <= x"00";
				WR_EN      <= '0';
				RD_EN      <= '0'; 
				CS         <= '0';
				ADD        <= std_logic_vector(to_unsigned(address, ADD'length));
        end case;    	
end process;	

End architecture;

