`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qWFZrf4WlrdSICSrvuOk4zvKVDeECzQSF4pssB4zvz83Pj/QQZEPv+rzQTslS1tg
TnSl5HAbQwNc+Mqu53tfTgWFDg2iUjWpg+CmAssojeCequ20O5ouZ+Y/nllk7BxP
h+u7+/FbB5tZHF5ORFhBr1RzwuINmRuHhfzPzkNYMohtlt9+dzJ974k09jmORSHG
n6l9rDPXO2/CB/xrFjbSRfJK4z+qv+y66iQOLazSpXlxamc1CwCnrMEAj1GVr/f/
vHZSAjrQBLBhAEOwikuSWk59VNjXT/YvFOP/ZIRbKsE4fbwlVzp2qVjSGsqTG7s5
iOvIn9/mNAvUeM5lYeDMYbi4NdPvgUgQEb+FUyrbcRX2MCv5Wtvsn6VljbsXclhH
ItByUnnGrOYVECUMWyyHQ4ECEPz43FGylIeaUNaLISliNBjkiLGizVaWloEKYG7I
aCE21T8aN8sHkIXpVLIV6Ma2sK17NhPmZuPhkv1vPHmYGr8edW0ds8Bw/CJkN3xq
+EYw5YSPex0Em/CKEX3c08HKtgtxSoV+d1oFlctcB2dgs/ciXt2v0kROnZa2v3AF
3mhsACL9xjQn6HKX0hC4SnWXVOU7PaybVcFqt9WsOXIdNAD9JPGcD4dXge7NfLQk
zMksE43Ud4WBM5e2Ksb1PA==
`protect END_PROTECTED
