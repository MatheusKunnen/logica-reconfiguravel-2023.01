`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dnyFboYdytn5Lq6vJtSK9d0chNMr/wConrRt6oS2s5OHT6zCpbAzHEWVWsGR8gM5
CRGSe5ZcUHatxceI6t+fUvfcQRh3yfGIe7kJGWZwGqz5V4P1s/dYTRegWlU2GdBx
YkWWj/bhRkYyNOJIH8tPfXYTaXWh0zoB13LP9MI6itMBG5RNajSkUenI1Wj4Ch1M
FddbcQWXa6GJjJnVKh8f1h9YU/OIameSVxtLfx5x3o4InVeFw2cyiSOaNiN/qKQv
eVh0bAcqlHM7N1GYwXs56wRAqQj6hFONsYSqpgzgIPF+s5TD9QFBHtZouXTt/wfA
rcTSzli+jThAyW2+HRS0Y2YWS8gFMrnXwDPkCYCerYbCpI9wROSAKA0jOD74GW6s
aGJBNhGMwEiipuwdkYyhoIL04YG9KiRmFU3kHJw1zy0AocXId9Wg00TK+1xpPYGS
09w2KOnR3dQaB3sV339EWsfn7VNX5XJpslrrqiKgvtEfM09nwwYgLhR4fU8TiL/w
lKatdobLov7mY0Nx+qy86cIUJHA2YFOU5DE1x03bFnTs9HW3nwNc6FzazOnZrdEw
H/ibSVDjjXMeuoAITvYSMGqGoA/FetfhoBykEEf95Ednu86Jv6s3o3ESIOxvvv0S
r7g/F72Fz5hA6A8Ul9bBHnGYsLPUF5YUJ8PO7rUhUDL7k/09p3cfPvM/RIWPduCz
1VScN2KxH40Q0weiJcLH9foXyWC3tMbgS2VgjE+pleWuks7ZSN6+7KebrLoBEq+S
oOK9+ZrRxHKz90NA2RrSXFhpXcneNgFgqcQuIgo32dzY85TUKy7agNoIbGEJS4RT
/eY4XBsSVOeeZ/fpaTa0LTcsrEtqNMVChSF3XQCV1zW3Lhum2DbbY551PwWty/Qk
T1enrX//aFTJEQD9Qxgz53wbK/uRVBQQOiiX2EtbMGafUWnZrs0cX5TESFTI/DIO
ynS9oj8D/kM3Gf8NNXPOGcTJfvQv2UN3tXHQzhIfWj/SlsqOs/MiHI/U8NGYoN7I
AArXl+rrAX5NCbYhQJNDK4UR4u6HKk/vfe1uRjeMT9bPo5qeOhlG+opvMfmxbkUS
pejGTFa5R5YmuLV2NKvVS0LzFeftJAXsxziTMFv8gA6MY1K58XToUHUdYxgkc0iT
bUjffpvlfaAj25NxKLKeoBnK8VCLJnXHfsNKc2Frfm9bbWJ0Iw+USI4L7t4tWv5N
JEsYDb7axKnUTeoapiCfvbfiJiXD1CaiDI6pk3zlnSSJ0Sr72jzi9u+2D8WDOkXm
FO3h80zFsUD+wLeaxijHmqRX3sqhNoLOrx0LSD5BZMsrKnt3sRXTr4jCL8VdSpUy
XVrGSwJjZwvC9OTpOaXuUPQe5IPFv0FtZtMnJUR7QWW4LEfQHDDQRRPgwyUHntNQ
UCP29SW7zSjGrl/Mvp1ds6lgeXvY2OSv/0+ldk+8sUiEwh6R01pcVOZRE4xgaR8R
pYzMD7u2Xjc3f6CqFyDLDiFhjycKXzsiVaqX+tTSb/9wm0ACj9ps7jWJz/nHlQFF
mOSse+GwnkEkYBOw7Ud8a054nbMdmmAhgWBQ3iDcpUKyO+6rvll2DJ6pZ268a208
BxNVYChcZkx/X2id4VydF6CaxeJwLSyD5ISB2ST7YcX/R7Bu2E0hIM0/lUGim2HE
LWuv7Aq1fRctAYU/h0In9SNnMvULlwUUchHS4syaeQX6RhPV+8qGGr1gbgIEZcUF
3HvUKwo7rdqMjHSLe4xVuAUCrLE1CdpH3CGOKCLGBZH70YqDr1Tj510MhqmtVN3H
8Ti5u9gdSQ33ymAVZMpNjk6sy27tNjp7oXMMngDAsGIkULXe7c8D9whAB+uqLOEG
Cft2rWZDR3CnrsafGTi/cMMnEhOkm5MLn6iKPCuVUlRXiAKmVRjcIlrmb045+8zf
xgdVkLjYxGxxlKD6tCat+CTtkv8L9mTKIMTgoVWgy1uZ2agcxA+H7A9k5obWK9YG
bh0ErhENnusdZHe4XyMXDt+FoCv5YlLwnp/gJxthBlqY520Q2xTv9sIygZKmaJYJ
/9rdqdP+qEIc/V1fD1uYCQOKZbPHaTE+2WGx10e/oB6YmbkQP+auD3lmOQCgo5LW
e4RK7H6XseVUjnBMF55DaGx2xTk2vj3GIEQSLe4n2OZZP+10jCHRvyYppJ/2657a
6XBHyxlhh/pLYGQc6JcOT+QGPterk2iIunFV+0Yuzt/M3DokbTozLjfmbTp59LDP
43rnVR2sKG1iLHAdb459LAlm4VoxdkicLeIln6WqL5aXypx319OsAixSS6NxCOVT
f4PkI3oBwYw++pL1rbI3CxRNytz8wc1ncg56J9IRa6pQD4H+cJy7Hzf7JixNK6kZ
NEINjBDODrKjXFh79e80wdqcp7xRS3EWOlZuiebcjM7O48HulDaPX/PZitsIS5/D
rkSpI/3Pxl30AmVzrlCuAvSaDz/Rj3kGLQNnt/xKNUEqspN2L1gl4Pr5y2h6zSXI
xwWn90vnv9Pa80i16P7qc+m/TFEeLrng1rvrz1XvqfNxowg1cbJFe+ZAaW3kgJ8i
zC5aliBX7haoaiBZB72nbHHHWaRZQ/iwk9Ng4HjO/pgPmmtMLRSzoptKC/EVmEj1
AfoQkfkyJLaW0mrlVkJ0LX29YOcfkT7V/BFjKHSdlJWdhmrmAApgKUnV28LStSlq
j682Zg0tcADKY3dcN2aNxMa24ysjpQJkpn/rVlMoeS2XPfgmNJdcFf1eFxZOs+89
x/nMi+ppYL3CGIo3JgT+Y/wWBrZUVGAyNoJGIaq6nvvUnP3gxcuEdlNmczmTEuDb
rDfkH6sNsLp5GdfqUlxga5Cp5Q74jzU6bpq6ansmkK8i+knGNTZi2R76ZksA7oaG
L6iu93MQ9BqhqrhGfMgVa/JlgBbXsvK0K4yoH3eTXlzE+gKHxI1Cek2kU+dR6Ppc
c0aTCKilBFwmwokASUzPYhOKjwq4BDuAO4LCArceXwfwMN92SFMIwZl4or8JCxsN
IL9v30V64DBHBwTSU6dgeTHgOnPp1jTvEE7kwIYQu3amthp87c0ZptVCNQg9bd5X
7gWEq5uGXq9xuwY9UBI9px6pJp5VR9QJmJLyhXsLIYsnBe201svkymKF2Y5aVfj7
gLunWqVXjfY9MZGJDYxDzEndR15aiQa2xoGE8AaLWOfcEmifWaQFiqo0n/72T1YP
JHaKyCwG+10moftJHJrak2xpB8lv5nSt2TTjfi8cZ4ZL3fI8KePNPrWAdaAMD2n1
qbf/zK6g7+aglt+HYhYaxSpbDQs+CA5utUmmYSX97MMCHBF4/tuOSwu7Q4GkbjCj
aFNOvwWhr6VAgy9VcMxNtIH5Eeic1MkO4W40dLgwjw0+5t55dveDSlHR1speuSIt
BWXULthhCyYKRyap1B6gk4pfUFGq724RZ3LhCbJzN/AJX62t61TFa6VkQ5/C2T1f
RJLYzkv21Hf2SoNbRKpc3rSv+90Qn/4zHeJ7Mx/Vbi7/WQpIZODWS475pxUUqC0x
eY5jk7zGZo/gPO4+mRPWrfLL4VuyTMXht0/S3oofv/z95ZdGvMe6TvW8txtn/LXl
VkSIuRrYV7bdD0HhfY+GKN5EiCQCHfpvN+eGHvMy/1DwqFmDlUb3Tw5V7swP8HAv
sVNwF9GeTgNbVuBu44AIMHfB54YRcBxh3TP7ESc/NElLw8xYw1w1zIpw+1UdesUs
Rj2cSPQrMckxhQjH088nq2lITFqNtyOCSr+yBBXSsKGV2PwHnxZNEpHL0L0dSLDm
8eEv1WUP8JLlPg/hWbf4mN3O4wGBCgdC1jLOPI+60c8XKJQ7usbpZlDKTrNlhIUR
nfWnNyB0zHlFGwfkSrMeM+z3XHiS4HXjrF9hRpdbgamXZRt74hyg/nRBg/Xrx/SG
Rtpb5AqjZ0psosyu++pm5RmdY7yQVqLwfgXia/4okMoKqFROwdx37IKGmTqsB7XW
wDKfwnwlbs22ulNZYTd3mYrtic3ogKlFLwSzQGQLCr2fHU5lLQXLBai1RfwhVTlV
i/0umxXTLDdEr3Su5UxaQOmnpcwcf45agTR/SNTpZI+Rxhpt1PSiP+Uj0328IotC
zRghqH1IbsEf6u2KuF7yGZDxk0yf8ClEOOOacTnARAoYniJ2i1MarJWx1ruktQvi
PJlJlzy1y0gyGHShWSNL86iMl69SLop5ADdCAzV7hOe70WQ9r3A/oeLy8gHNB/fr
HE5sD7bm2aY/sbhykHbNjPIEeUgdJFiqHLRYHAy5lc7j5rS32H0OKFNvi8XgeXO2
ltAFf+/jKzhEEE1be6xrtxTnjvVC7rwPV7bgiQu4bKpTHZIxHSL6ISRp2YvVgWow
qf1ucWZu50Zu4B7YaWJ0QizmufMRiCVltf24uV/BiwaLp3XZbdRvACjbCA+RKR/J
GZglwl7OseMf+hSejh4JOSGAh8wG6rX32dPZqENViTu9UedjJr3s9Adf8LZYJIWf
AurxCePG7ohusXhypulJTXWe/oI9ooI+eaK4sw0P3eCKRBfklZvVGa3/8OtGUDFW
SKUcT6x/hq4KdSEHsdLe8mFGXZgvEB7zpjzgzTTVgmwnzWxaucuQnFCSZVJyVjIG
oFuAgZ4TBCjZaMy2uAKXbfxQSq7gkEObQoYy9W7x2VfMvnDKG12tQn9Xz/BZu/Dy
lOaFX2LW5aP7XbCArs2We9HsomnFsIYrUNqYNWIFpIs64+g7QlVZtz8na/LS08w6
eTZgnHffMyWe+OzhKc23Lfnfvm66b1/YrbtYGxeM4hL8BLfGsKdvTsq/g9HZa3S2
UiqXvBuj5IB0V0+MNX3PATlJi3AnuCY11Xz4X7clkqk759LW1PZdlRRJEenPvptP
EsCA9eUu1vEtojyT7j7aWEPkdTuIIJ+nVAJmhqRDD+N5IU505AQiExCh6SY8eUmO
pDceqBb+jnF3C6hH00/poWcGokJDU6s7NisIGz4gKpN9qNZJy6f9qcwHWr52WtIg
vkdPuXFe/TcSC4B+dQiKnlC88XFqiW5ykpOrqKhPIqhOsueZm5WnPsxjglBrMi1N
khoScSdPR/DlpeJTYZBl27ZNbyozH4nC6EBTl0UYDFdJBPmh0eXIlGvyI3S5I9vG
YWbSSWqo5IhAqvDnCZ61tA0BBcYf7BZPaTYqhv0ChL1YRy1nCh0J5uoLAs+31x12
8G8pDPlQS5Mmjzq4RGE2z6T7d1YLvfUgBR7dwP2M1ALJh2ZikpcBsyPs4eThSn8z
IH0xL8wFLFybBGJsYW7D9p9itIyAvgXOXD4QtN4BHF2gSL1S+hA7ABCRB5rp/GWM
lS4j/PUUu0VJbz2PCJG1T1kHv9btVoGnrml8kLMlpY6ZwbbPzB/2THxgwEzoGWiv
sXcbd7FtahIdcSrMmZZcadP8pMTst8iLn8s+eobtfLvLsXXDhW+ZypWxqOqvNFzV
l/pncmInNiv4i1Hr6xm0w04PuqgRdRfYO8Ch9WdQDScczLI9NblrRhXPr1zEIHUx
5oB12Q//jEgn4ToKurkbym0dJNJw1dfhFa7MovlTorYzcwSOu2erQuO9PbXRPrKM
j3joCGibDEqcBNIcqz0muN7ofUmEApS8KJvxY9/1+pE73sZ7OFvkLqZ+/7i6vPvY
NBYd/kpQm9yiEpc3GVi19cxPBm1QJLBa+DI3mRw5rW/OVWiMAIc1+J7otwXefCl+
kmF2Jihwbrq+k6YjUX0r0ykjagvmOzNoGCSxc/sqnwYOXDV+IMhXBWDBkDZ0s3Wp
+sur3ENLH7gw5GyS3OfCerMbrMwpoykGZv3ldMVymZ/EnFPwswC0KpXN7YQmAg3s
itKR0Mi8A/tnp1ktwCoRZScO8dIHy68bSS2+oxtodJ4ValWsCkxkSfBbFzm3Ryhv
tZQ+pBv07Avmm4TNQBNxVpIdYv+lqMyB7X5yGQwnZR424nZ97P889QtWlLwTm9nF
DnCSuiNagFyaBBOG66purTeOZHBQ5thD80RekT937p0DNYT5Xk6YLTscWvx0y2vA
v31clcQEUT0NRE0bjhcK1iXZzo0qpE7jMx+JiZW8q/0oUlQ78gUjGKPeM/KN5HGX
Sh/OWEYA3+XJHP8PQ8XdRIBEw03bwWa4WRbNsxsvvq1ClK6Jl7JS4USQg4N0hFbV
I+iWz8xn9wTauCKd4IrvUL/K7UdtqToGK4MxtNmcvbDBz0W2iAbydFgG6N/m6zVk
q00AnvG+eHGkjKIdm3sZBzh5bOX3Fxy5OQzFiw9JpDLhPp/UGePeMrWTVbSRC4BY
0sBqgHJX/grFYHWZFE1RUoj+LHobTu80h/x2WSuV+PPkDKKyaDXkidqDgUiuiI/4
Pg3lI0fuBfXn9yL7wcYmWnQTk2EezBnVpP0dXU5RVQxDsxW0HtNPeR2xGI6dE55Z
ZMzZdv2J26MKe1JJL9dkD6I2yl89sbyxHsj1RhhyPzu1QY8/TSzELZfOapDuPcTq
jWBsc9oJdLK0bjaAqldvWm2YpeKN4Zz+Pl+ByVHczSADNctkm5KQp35hN6dfsPpq
SjnRgPKaInf1C0wmMsvoJvza38vkbLDU/dC2oYcI8EXcygB4t2m44TmoRY8iikNh
9VvCPP9644aSEbQQd9djoEDXr/DgX9ZvYsZx7ksf3+s0sXuSJ6qPAbBMDRASta/6
8p+rFT5J8g65SjyfBE6EMuu933kKNy4lRXIIpQegqGoLaM9pvUSC5b4BW1GPasSy
sDSQVb4wU3i8Ed73CS6d5NFBHIsISMOL3nAVPED9kZaP0fhUWWg+v5zC/k7HkDi+
ntUIPbPlphYw8MFmG/IopRIHYA4hjK11BPn3Bhe/cxKkwNjzv4VCVSOmPKb6lMfg
sQa7xi4iVnqt2c1xxZVDYVq8Oh/rfAhhN6cv+jmWHQ0XO67VT2IxDNjhVGO943n6
krETUAsw02d0MQBvsng1f5cDbJU8arup9QE6wPVN+HC/pQx6zjO+lcZJ8gJ219HZ
ZuYeeLJpI7CB2aMMHM+1IxDbOvEPJSgE3PIA3u7usORSv7ep8WDBgFULPyzQJflJ
fJ2/6u+fp7rhLLibX0dpUwSIeHIZYnrhFcc+REzJV4Irq5Sx3/gSjATCr0/vwkU7
Z95Q0dY+25AuXXu0bshjJMGqfdRTQaptdrE9qZMiDgVXxL44WLeTJY17ZpRSjK0V
UnhiKqK2Tz8gT64kh98KkO/mtd+tl3yFYS+faLpl2AFu/rLeCEX7PicrxMPjsZuO
TDQq91lkRWrOe3UKzbhsXgMnCLTR1ZD+OnJ3pyFv3CLo3hxUREe+RJ1Lc9hvwS6e
V1u+ViB+qYFp/5PHxbZ0S9RVoSctXCUnY1c7BBODrhB/MaReMyF+CCU5bVF6AWBc
6WfP5kXRUT8k43n08mzgGr+RgNjCNBVi/ZEqnMopDR71iUtp9zVypUgyNDFFJlgq
6WNHHqFj0logZSatBvJcKbZVBVKmJWDvF8Y8/8aFiKcoUY4KhO0d34/V2UlsIzK0
jv9Y31R7k31TPsCvXj1+adctX9HbDGbZybk+nVQ+KPT2V24qjou/95EIMAuY924s
Hf408ITaHkkJy6uo79DwPLUtcja2weqJjb2uGPGnBYvdtVTT8R+F3+BcVUTstM0k
MT2CH0h6BLvS17m/HQznWplN1eeM4TDgddeqc33PqQzdf2AIWrXqrknCdZP4cS7O
YaYvty/Es2Y1LUiK6PIT5BKvTC9jX5p/LlJtn+L1j2W/TN8ERAMmjeNlxp63xCMl
MMcNfpVR18Mpy11mp6MVSprY/J8fcWjgLAknT313DdA8DBdU+OKElh1V5/NuKOv0
3Evhi/ZW/Vy+ZwShHC0GSsNTloZv1qZMHZLXsiTT1k7KyvZOaD4DSM18dP08oxXl
PDT1jbeukgAcQ3aMn9djHqAYJNRhUqnTdZPVk/UfBWByWe8nrjwetCGNFB8Wl8ZZ
8TitWkK9u+1sRzfF2XMQmmB5AryzukNTJjmERkTLTbx1+AmbQPs3zGRZwi+J2o8T
fnd500mKdV4d9W8mJ0KqsTalc8zVj1wamYgXrtzEcNcic9PbLQ2tV3KXoyPo98Mw
cZ9QEtho5iU92GK/CuMRwpY+kcMdycWYyMMdZk91mKusOBCtnzC/lhoaXQnD7t7x
qFyhGWL08QxO+tFUIp4xMIlN5qfav1LmtK7jtCbpgbIIGwWDKauUP3LMZqHlugYv
Hwsv1t6T+ew4zb2EHRCmZzznfg0GWMZhYbQzHF5rHO8Q0UI8CV9fccGkuc8yP2tL
IK71CpdwScaSQOax5mq5P3QeSDI8BdZThhLmufy0ubvYggSGUwRrFdypaODivAUV
e/g1RsHVFkgIIM3lAi4umdTcVM4wXPyyUFhwv2ihVBgdiCE1UGP/0oeAnLKYdkYr
uC2RQOPDzGhTtHBOpepYoQpU5IJ3TncBc8sVmZ7ManDHsoxPvRwneQr6+g1z5BzG
v44YTKtN27x/3so4TCFTJ3p3DGJF0EQwhbiwlXvsSIShBqgpCgIjjv0IatywpZsH
98a6DiB0q/4zkSBeo+UUTy25UYh2J+u+3KG7SF7ctTmAKLXZCrKZ5914HEtRwXnp
vy902g7TH/LmVmFXqNegZdyq9K+6ZADZ7qFqb7Fjlhia8iF+zm/hYhVfOV6hr2cK
+o4yLivTE8/zoqtzsPjuYB4UpW5MTR9hrPOE8cTXijVAtWb2k9iAkz+oCNFiMsto
59NsLopDcqbr+HWkJnCgdOw9ll3KBWrZNbF/KduC5B85i3Bxo7IELCCFoP7WFtxM
RzgTHOClEF4VKWm4kF0bn3lT4xSKQfMX3HVmsLLwk5APtwEBcB0j52c94Y2EyTy5
fte5+D74T02pyRZCrp8Zd4UlY0xY5z19SkHYy1+x6Q1HI0Po8CIxe1rNaIoBvKOJ
/cIMD6/kebxqys8s4va7GfRsihMvw5m8Yhax56SpRyw=
`protect END_PROTECTED
