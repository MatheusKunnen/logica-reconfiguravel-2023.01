`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
onbb6I78zguiLrE2QwOWnaB4DYE2aXXD+o7MImXlE5BvrDHKCAYQXSi5JYR9NDga
Rxm6LfcVj+8MuYiaB2gitLNS+IvzNOwB8Yf/ObPwgjZRSTUhDfsC8oaFFK+CKVki
RXlNFHBbG6JCFc0a2VcgTq4eGFChgtDnTY5JBqomWhUt8EGl528IQS6bgCsqLUNZ
GVG8aosx4PitPz5hA+qzzvamk2OSx6LEOFmeC0B/o2lqKAuDqzDxfyQb6Y8ExxLQ
LNIgtgzvdQN/ljIxHKIqYxvJY/nuS24PHKPEZ6j2LomcEF/xo7CIRZ5XOFdS8IOW
OiuJsYmoF503hwmSiOE9lCm7EjqoK+rWhBUwlyITOsQGLoWEalSRT2SnBVG2jyhm
2DGNFMgcWfp9kqPKevkN1Kz7szC85Ncr58QdoNCHqEPyQPaXPjvKXZH1NIr99/C5
atqNzKkpOMTe/Y66ksQ+od8F3qrT5YHhj4ZZD/pIFFP9+fHcU68JlJSbIMc+V7ef
xav3kXJ51PzCiZdf7phf4UsR8gII60k+dNziqD9ikCC1TzWx7kqkRgTnyzMJFOQ5
XG+b/ln4jADqgUc7BJA8XJDjgnS/PaG0+Rz4eXaaRESK0P223g0+PZ2dXNl4gVdn
Jx4V9+XrSOs4DhWdW0PFv1QEKSMXPbyTzvBMK38rhtIB9/2Hjdd3Mdjl0dpUzAmi
xbsy4+FyD03NjZEh1mOKPmnbVNzlzAHcheb5mrXcP0s=
`protect END_PROTECTED
