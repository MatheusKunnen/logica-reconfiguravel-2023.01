`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lsqtIP2DInWzMFgJx1DlSMZljJq24hBGWazvd8X1OzWIApLaj80oJn1NzVon/IIo
A7LEVP3onTczGQiuXPhINUEdOngduFdJSv7YOXfzN/FczltzMT8ko9oLVLWIcyUz
0qByw+NwUEOs8kgmBQWR3ZyM25rs1CgmZabAcMkuTZVXYSdTJaZlm9Yh6vhqyfV5
0P4s0bg2NxQJLHMlulbuVJNRfNX4U/ahFjoS8HrxEcZNUA7QNG1c9qVQGQzrClvF
7vLi0ZzuCtE/DErSHAIgyOL0vNSsEGjlqjrDrItYTVezrVULQS1/Nfrn+acS3cr6
0lgAwhC8DHgwfZAxbCGGTcKoojt5opXeZC8OAElZj8zNJCWMuhp1iABJeSgJxWjI
Q1J+SSM39UCi9SX7XlBB96/wvfWn3ol16ry6stjSh0jWLfMDWWBUVdkuiL+NXLMq
x/QqghfVpBTnO+LjYppOJjzujffHAxdBiLlewSsoC4d0ubdITsUWy4TaHMY5jvI2
D+N8avrGJaoIR5+Oh+7OuBZFvto7pyFDacLaJD9C7BEtvaRiKjm2FdBgn6EG8lj1
gAFsK+ks8I5a2uJS2Ka2tucWMCDK3kpGp1veRRt4frMIt9e/S6+XNNO0zXAjJ74p
Zbtgsgu5ee1nhmgioVcRnzJWpU6tiZ+Lf5kbK5vqquw/JdH5BKzhf5p5/YBqclPp
iQLmWMUy8L1IyzClEuAq1h6yTQwt6LbfS3ofHUtdRqovXAs1Zbila/RT1a9cEu1f
1+aK9FHnl24x5g/loh5wcSVhRpaQOoBwQ4XnJ30s2yoOmeQRiB/W1m1C/bKa3YHK
5TxgSYHgl5Ee5fkGquTgPAb5d2cKg8ehyMm7xouAPeNDeNpbhZkSpL0K9WjQv4RM
/X/BEoO7LJ7q44ZyV+8KnVhh/kKWhqJJuJJQ90mcuQyy0gD9sd4HLFXzV4n7sWgI
BVqhJn2sliEUlnT/0TA1a5r9ZV1XoHAACGtEZSL3UWLsFAEEWEjpHnXtMZteu475
ao35e0dHWbLd5v7FJ+umXaC9nuMzXPZzJDsG4IWQYDmmloFa2qOnwwVpp0tC/1OI
VAl1woJArt4kVo38cHMi6BoxWtjM+fzUxyb+6JOzmI2iYa76tkvwOfc8JMnml9lJ
q2Kw753DM5m9Em7iUWsykgSrrLop9QRJpMcEx+k6OET3MPxVMXze6N05rv8Kn3Wz
9BHywhvp14zH1bKOzNwBC9j+ZJO2+SxUXvHIS3Dk/LVsy8LmUmVPYu4C35LpRv0m
Zs84TkrJhwbi3vAF0lxaJjLAAboYP2TcmzdZEst5H3ltpk3aHY7ziFITP9SL5Ilr
4uNveq0mORjKMkaFQCnZo1kr/QXEK5G+t/MV+f3mYitGLe23KSwHrVsdbXahNJCp
4bfN27mzh3TZZH4BdpGjy9Cw/0NBOu1YoQg6ikSvUlbPNzV+boRbZuX9ATzB8EnI
e4PncFxJz5mDKKsRWCdakcZJphzta21VVD/xBfxRVfpLBM3SrTthRYjVoeKDPrbi
RLct5SpgC1A2ogm6sBFZ+YrLEx5OkywWG6hMo3JzthERoxwo+DIcSIu8lTTz0OMN
B+Fid6qQZH4XpETmeKqhCzDAyAY4EUsbiZ8sY+DcoRYO7gp6kvf43XEXrSWgA/ME
MX89lcONvzlKDR2xcUGURBX2SOq6chZvmFhM9Ca3kfwkyEERFIsqpJH28RwVaNIW
XmiXAYk8G2uNGUcsxVDvT/zNt0i7sY1iR33vl/RxynStGHv0fz2LMXiGNsNwB3aw
D+iNWf35rWYueeRBmopjBH032o8qkquge0oIiqtpOljKhpAdQDW4UFoR+fngDpkr
G2AOWIGmWbLuViOZ8gDIQ5hjpJOUmB3jhDXVIIZ51UX0NRd3NEsRKe6SAy8nx/7A
ExA8OdugdfZ02vOdMwE4JRr36Bl1XONZa5c4CnR6dqSFSqtoJX5Mm7Uc6nLIkTEt
cM0KblZb4cxmbWUGQ3DGG3gE8+yZu2OVO5eNp8mRMeGDgFGmoRfQjR1lnnaJe7LR
iOiZVLQuBGLut68wCNAoUEMGb+jq51mN2741m1qogassdrdu5H/p2gFLRZsobVgu
MuHVEnTVzGWLBq0rFcRXnb/hSjpIb0ZBKXhVpmwAw+0w2LPuNSxu1btpPdkcXxNW
tOSgpFNmJD4fZXn/AfJgEf/e1bpcJDQG9Bt+9DyKedwhJUgjtJEVSh29QVlb4XP6
kgA1HUe03MNPuIxKJ9bMng==
`protect END_PROTECTED
