`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LHx327Phv8Ety8InHPjA64I4uNNMyVk34vVDfm42sKS3JqDbIeXZmu5XtO/5Va32
c4glR6BFnonAs9mGiEiO6UD9mKs3V03G4aBmrw4Q7xyanu68oo/IaouA0lxchjU0
nDPuthRj6iK9xCRS+5inp76dQUXmGOq/FwWHO7c+iyDyBMprck6PN/EqxUNfrMdN
JzADYoa/bIh9G3JENRxedL55QaaudTwtjG9F3n63hjzkynEChBtarLXvhvy0vLhb
/WZWzPov8VelH9Lm+lrcOvmmJJgB102xgbGfzi1RClBywmSdcIpZ+eYQKIbVBOQT
AyA3+XcBW2AQp09VRUr7c/VGG77ugySkQfhQkUaTP6d7eUA0WAnA5NzPm11NKymg
xHK2FVJN/xyMLqSJSPPDxI39lkwVPqerIfONhM9mEZBH6p9PQ3aiHIeURV9r7kKb
A3VTUtfBDoAqm2Id6ZDEngniuslCCFbEKwYkQiK2jfo+CBUuFEQ/pOaHLREIzjgQ
5DDUQ0hv7IcMEDMmYFZ+egCFXwjEcuoxC4vl+OhlBDXQsYKms4uUkGjQNDrbDU0D
/oLFsuWUjQpI1wbF2JQaYQvU1XxzfqT4sVeIsxKEUnD2tyNY6p2or94luFROcuw/
tJQLV6XqXOTJN1m64T38eWbxlpWpDA2zXX/wYGfA3fadu8CGg8uI6H/BG6gIqsQC
oSx1to6Bn4OfmHi4t15Kcggb+AEQ/COt776UApgIcxMUNQ9SqQc5yIO0/3Zqa+2f
tb3Kb6N3GhKeUhp2fGWq3+skSSsxe51q5Az1glNCWZoHr4NGwfz/aYh/OsECITZO
qEo7pXYm+sdFr1mApB5x0xFkLefOCFqBjpb8/UTUUj8LS0k4vToS16/JaHmin+tY
SV+74ph9ltm8VeBqB/cgwQyYB+m6pPgrddYoi6dr9LAIBS/MELgOyceoa+Qz6xtQ
l6Hwb2r7PZS3y/Y09MEpL9fdnzrERNuvIzvM2/VfLF/czBvxGFUwkfMSg3fo9rx1
YdQC4BdHkGW14JUsjR4Mz/ftoB/JdasPuuSaLGHbyY1EuFG6IATI5s1xnKH5Zx9i
IcM12QiIMgGELBEyGVs6Lsq2e47TKWNmjUmnsYCP0Qlq/ChAfxPNG8aSpbuXtAe2
tPqnb1kt8RX+SCrTXjxcjuHdlyN7LbQj1HwyODR+KHHNon3z/mSsjUL6y6r0RYDg
GeVmbK8PVe+uMeWYHSffWi6oCiHZLNnQ3u6VG04nPzSlEjELHpo6XaX42wf5S1iv
8zKNq7T15DlAHNmpz4pZ439gczQm/AEsHaNxlIXZGyN7hdBEu+s4Ybz5RQccEhCI
S5lX30IIkYhT5W6Mcz3tDg8OwevsSsDl6avqg4Ge30p0y3DdRqyuM44mILjDnDLC
nrU8nposmX1w4cqGTs1wxne2t4sXyhn6zU60ZLAPN9QAIzmHj6OQ/Clue2kYMlws
RA72oXz60B+hF96jsekboDVNiFaHPwMEA7RdzznKBse4K95UqcNVRYYGM31QkLq/
qmHCVaq6PXMsP8nEAFNCnD95BCH8lUoJTxupcWyy35e3p7v4rtT2Ok3PxfAGp7yo
0FP+VFpgluZf3jmXWJau7cS1YzgV5eqL6D6f2nSHiUAhcAoF4hapHuomsLst5KPf
9OnxtNwhLu0W9VFVNqjXjqJRRovSd+xhAIEtp7uhFod9jnjIys78DCpB0lFpJFEF
SBQOjUb7jy9qrG55iHUjskjj4UgmqjEaxTKTlwTMr9/oRz4BjXcKU4JpPUoGDvQ4
mrHYWAlpf4bdF80uEBFT0Y4ksYegyZpXb+7yoBWOjxKB2yiQPO7dF33jns7Fowjd
B8DGD8bPYlE8T3sJca/0+UaEhnO/7tk92z91722om9/wDEUysqNvYrWYNTPWbDdR
GN++t7SF85XlEc2q2chWP1mI7tK38LcLRT2lBbGQoQnK9A5OveW0ARiJcFnXU3RT
LeOtLiLZ+Nbx4nIA+auB/hkeLDITupsNbMCYZUbxLAhOcJ/hsfpqv7tFjgMtCsYm
n44EEflbLoqziLotgmxelBcsdOnzXNSuj2pKuP25u2ehN/zdbNkii6YrOR4z5hOD
Dp4ROLYsjyXin/yCZ8uL8kw4/LkSh2kkSz1YiOGJ7OBo3Dgm9HXviiIhyvsI9h+E
EcdnGugEiU/td9TOHUeyopaC9A/Iec7jWxEe5xzQmM8zPapmQAgQOivBkWzFfV5P
QbgxwYpfCK92URefRAkeGPJb/W7ebakqTgLDnQz9GDuGBV2ENxwfLkvzw0b5ZMsg
njv467vy8nZD+DRe9wnIEby+8v05xRhouw87vlX+xnsFOIa3E2QGMx7/3DNwVho5
2H4d+UkXZokmXAwNdg5ShXaYzKLFLPztJjKCuOvMQ/4cQMyzRsxSDmXOcUlSuF8t
/+YTUURV2xn1a3vI4wlMPmy3Dnr/NoBYsTj7YNp+wKXj3ZRahu0QCWMUCb+eiUlz
T2bCiWkRYJOQytYlkFhvozDGyUXvBqqRaGJES2UPz8+pVTZ22lK6vlj9H5n+59u0
KMNPdSWfQlks9o0vLd2FsTyGoWkclq5+G4CqBqQqQKUFaMcjgE+PDZhELlXN8Q4z
NXS3dnzK8tsInlMhqBqVn4Ga60bRxhwnWB2xgr3UHzyV6ZJZxn0Q1DTySCfOUJop
biZuAP6ngWEB+hIFi+ZO6j5tefsBJN7xBz1n9SFIvyeHTscEKSSFjagJJJaI9bat
+++A8qTXO0m0q+TG9h+3FmPQDwz1NVt+ALUQb2+/5pQNc9BgT26Xp4HUMYnB+35U
1KqP7HFga5zBbBtj0xuf+F1+r4ZVVCOhjDNbekomIuBxuvrwsB5UgWV+vGIVJWKe
lkCFA1r8ZAB8xnhbscsLgJxUn957lYNrKdV+4menbOhCL7DzoVpMz2/NsO3cAND2
pFQ3YPu16VFRrO36HteeH8MJnKwnX3gMfnDEmUBNpMsc4LDt7mMDeX5rgmBBCt8i
nD2WqEsZKYgRTMG3UD68zk0SOLADEABQ/Uro9paE88+pwAYasFXZDtjqt/8M8jgR
he7x2sd1ZWpI2RuqVmItzDTHm6BcerWt+VAVwmPfUdZ9THQWO0eRPotomh2zEl4R
nm+ApAeKZoQ80U/RLP0gY42Ytf0Z3uh1hRZKDhhAjfRZboXmuURJ0Xg78jha1E0p
5pH7nXF8XOB15z06cdWCBAg8myDVJeDN5XlunDk1fTt3Z3qqyLTszEuitwj3hJyv
xu+IQpceUTaPgPElttCGQFfcddgCkWR8lXBL9bz6o32/MJiFuaQcqZZbAfLJdtWA
EFtuqI2pQFYdPCG31WhWQs5NtvNISPNS9Gty1oVGFIUzl1EPXwVgt7x6IWfbs2L4
9eK13vmg4tdVoQvyeCOes+j+dxaVGNH6DEC7bVTtYV3zF1+N0chEgz/fgxDqQmtD
t7SoV67d3UiZrW8hSFDkmYjCv/G0mPC0mXGW4/KeS92NAiv7ab/HHJjA8Xl32vXb
q2zelDipGWtHty0zqwIChi1Bdv//zLcaW7z7YF2M6PYTKWCgMrj2kxdyifP1Ngh4
sa94yExVfrSvbJLiVKZrRDdBG/mORG3b6gfcCXCH1D1dEgoGvpSv6ADnHACAr5Ja
yv8deC+OdGEdLuZGewy4o3sBE23+lGF6m0AB61WDX+vDN/rILCG/TCp802m4N9Dy
OW8+tbLdp3ehDAzOoNZQ8/Ip2Ee71rpe/bqKvLRqulxP0dk5HYpKtuHBObKhe//v
muxWShmbEOROCyFhtuHZuRo0tye7KhGtoIDFLsBeKyKgvri7w88Vpq+KQf3nN5UZ
5PKH2gy+hem9pRsyVr7CpRq54KSIEv3OYzaFjIahtKOisFopqhZg/9hFMXdF5kUn
Pkb2OS6pYsVxA3lVirclPXMhSo63cjlwdK6Mpi8TohtoikCqsN9WhbzbLQ4T5lSJ
1EPtwwdvf/+tjNvML1+He0xdJF5cGIzfsbM9je7RE2r5bQpJgswGTpO3pM2ChLPk
Lf0DgVQ5akoGHCueJCWdWlw+Hbgdf0evasswzj84aBXjL/zL5QEfpHYDqx0zAT7j
wSoGVAjTF4x5Y+t3AXCDATVI93B7mb3Wu/Yl8iYIWo0Aa7l6IO5btG2akcGvPfMc
8szEc3voDx1ijdOai/9LSvZ6QH/EqkN84f9di58iHldex87VFh1jMsnZrvl/mm+r
RdSkLkk+iSf5UzcXQu7i9mchMSCAFtnUXOD4GKuQaO49ZRPIk/44pMNBrYcmAvcm
R0kZxIjajcaB9x72YlrKkFiPxKl+kso4rDQUHjbVHUtNJyci5iA54Rt4r9jRRKj5
WJ9MvXFxcNBZJzCDp+af1mRP78g6M0orqUmcwZgKRaa7yOHpLNLkbOcRz96C0gMM
ToG0or/8vPxZgqt7ftK9hjOYUml0cRpoEzrUqPZKixZNbATIw6ShwwBoJqUEFSww
nfeW90BLzkJ7H4CGqwvrBFPzwwN6TeBLJr5Gai5EXECf9IxFWc/Anp62objjW9DT
nvHm5lrw2CwC4uM8rmLJ9CM8yTlx2rbjY/foozA9UZnlkmnliyVx80m3VC8/9A/F
WGlepTJ6eNIZivj2aiKBlIzKFXaeBw3yWiyqdR3N0vpZpImPUiiel4zNYlT97mdP
BAuP1eIQfQ+TbOaNSQgXu4Nfb9Z7kZvdKa93+AClGzBATdl/0ivj+8j8Q7Remmim
aQLP7nNl4/D6wTdc6s8bcSxLVaZyVi2HT/NigZ6BaiPKFs2hL3EaaIZcweOA1JiV
jhbPi/ApSTaR978s3y75NPgVIylhSVBcUcDvEwZLrX70z07TiomPGZbK8DQx3RQf
V7/oRlsol7qLAXIVKxMs8UzHc84p9Ba03gT25tahVPTxU8v1W7JdAIY11vDdLNyg
g35EEvsQDuQM3/l6sksFTB5K4Bnldomb1JCa2i0FZteR0jec5DMuRw0W1J9n+7E8
EHZdyL1fKVJ2KzGsYCHTO0QpE2UExXjg5GoRNPwupOalfhDW/9QUmlY8bkv0opG8
wrqN2HDBWhIE9z7udakqpJh263bdPBjttcgisy+qizo6mv8fSnpnT/smMV82Mu/e
KuerGhvb5aJpyzooOoEeGYlk49QT3WTUHDMqSHyTGsQQr2VlUtJIIAGKa1fSxEks
KmbfhK5LG4l4YNRFgu8mMlouUx9WqyM+IQi9YGluCsFulBVHmo/a54tRLQOyH1Z7
TrEz8LRyzTdrD7WNLZu01M1ctkTNW527xBwSBDNEj2v9j8vKnu/EpqK6//ab2JDl
jdp/AlOxkij3Fbh55cEyQG0HcjKI9QcQCVwJ4UZc0zlVS8ai3nDY9teA4k7dEVB9
Hp7HppV3qsrjRVEG/qDNifX+n5V5vKNrGDEcwozXvQtCYUenuEeIsMKTq946MeEi
cGgW0HGTt5jzLZFr5Kmv0T+QqDEFzWv+PF+Dn06Mp5fYVNeeaEbtcJImrMw4WpRs
3CivqyS49LUIX6Srmoaub9eN9zW22d+QElTj73kfzf1gUY8mV5gjWUfzIUI7O02s
HmFTMbS7U87GwmFzLCmnDfFlQRchnmKuqowHQzoLOnJQi/b+BsOnOgP1eGdWpnJh
JPAI007qQYeies3cHWYaDgjTYyTSdY89lBKIEpGrw4Wbfb9oHN72TqG3S6jmmL22
xv/w/tC3WC/XCAyT9CJfRAISv1MUr9pY8C0H2gahrU9QOBe/V+PmSbHw6EYwElxN
+cIJE+MpLXe5gD81vpwrV0dzLTYFjpvHVCJaAssVQxmL3y3rxqlDZ/UiuGNK7Zfr
jKdxtm5ROP27mTAeqRDBWD0fkw3maXUNkVWWB0iK4mhtIOeDjfU0BfIpbQyVPukt
P94kWVIcOM7Zqsn/2YDbQqnyoFsASJPoHk0D36/4HfoG1TN832AL6BHijDNoPdsN
KbYvxtiGHr2prT7q7vVvTHIW8+PicgCM0SLw4rs0cpyaAmLu15gfQVutfOZ4qOJ5
g1ZU32435wHehMjwA4EXcJJ+7NlB+FZV/XBOY0y7jvfVwfKUGflnA0NkkL0CyCzV
/Ur5xhPKuKK2bjsDqfdWXgVgraWG4ib1mMGc/WMy9m9nYrWg/gJfV2qVIhkLn4mO
Yuoql5XaOQur5j5IyTbPjO7Uxxy3f2Fv0Y/CMbv41zN855rZXu9Q27tHutYaDKym
7npzGwnL/X6k7/tOAxYYe+MUzvSaklL5yCWyKbU2uKY09TxTCFkKCNH/bFkqAIrY
i0G461uim80183poqkxh3Y/E62KHLLy/S4b9gubL9DXHk5IAqNj8nW4D0bDjKgzb
X95K3yg/TuerX/cpBMgRGCoeup69pLHBrBVV06/VrgBhrTF2mfVA0lPtBWywL1D3
jWfGrZmf419q1cyPF4o6b5CCBBeQeWtiZqsg4Vgairu5h0PkyxFJ7oc8kQgfoh8w
zs1/CPXYTcl9GzDMLwzUYWRKrihPmck/5xjOGWSAfytoGwJ7c1PfQuAN3gQXYtJu
RqASjfp4nMuMIB2BtnNendpjmJDK3Orugt+2Z7iXhS9jF05XsSamVsZT2JjzZlTm
KHoA441nYaGnACDx4slJJZ0wNFssJJaxMuKupIcKCZyMcHAJG/cxzXbsxxTOTJYu
2T3ZCP9oO2Rhbpk81TcJadY7zIP87wB3KqFlFjcBFik=
`protect END_PROTECTED
