`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wezxhqHIVx+vW4zB740RLPPnkvzNSqXn7/ZteflXbNaFkrX6DtUKRs8J3n8mUjJO
xcpQpNShQ94QtPwSXOosJKDAVowyLeTP1srFsDNvkPemNYhODgTYs4M4uwdoaRpj
03arFsjywvkka10zng3gbvpJFt7U5Wmc6I9hsHIXnfDO7EIJbbcU4D4IwUUizqeI
uQwthbagI2/hFIOi58nXhlQPFYf/8HOIeTxFmmK3Ym7crBvrQ70IYdNfmiuaY1Ls
LtwcwsBSchAFOklIN8i4RzTaJ1J4sNz8e/R1rERbk+eVYlTOG8N6QqoVDBS6DPM+
sjPNWDsq3B0vCVaSWudLmvHdoSft+o4XEBIK8ZPjgyO/Wl6/4rFwKrHnO78QHBbg
fM32H3H8mso3s/Ptnjy0NyWgcRfJdWDuDf9AfVRRY74GD2ee3ZNZw3843nrqXFqE
Gs52oZ/cs2oS+XMnsuNRZTO06Xr31VAw7FC5yZG5ZPPacXEMQkNjqEbxAHSQrxyq
ZsSv20MZvhkBSBA8r7TkvOevXUE7yQP7FPrepTFuO4lYRvdJoZjq5cC/d2T/d/Js
CSZ6cg2PG0fGyg4EwKK6FAlx3psVkaso6NcpDrkFCqvqgPvpv4N35K7WF4oS4Jif
zl4yEhhR0fI0kjKoSmv40e3zbc4d2u28QiIKJNbsEwfxkFPpiiblRvBdQMm2A2tQ
unVuqNlOgrHB9PQJTWuv1VziELyvl1Bp+hL9Sbll+qlVOLeTSwBiTe3QfOR4RnQO
4jlp9ChYHSh+7cyZGpkaoweh3B/WVSZwjDyg5RH5Ktil6XsbzKMg0zozfYy19i4q
Q1sbtL9YWh8z2wPtKcDTW8MJ//2/a//tV0fsS2ifYwVvgLzxC2Q3VuMRgXumsN9I
tFvncziSc8CY88Lkl7OM8j5hsXoaGsaQ7OpLHZN2upab2qW/0LR/GSsm5IzhgK8U
B5FXs8LeUnLmQpRY2ANbDza7xXpEbAtnOnIBmQsVzjY/JgL+e1IH/l2znzXv9GEF
Eb23amRQmeKEaZHgkI9XdPaaYIOzUX5ZYpCobHBzWcpew7z02HsezRa4Gkfrd+lP
DlRhab6iJO2e5/Isadc/1JDMWZs5Bg8q8VpD7M48iRIKRs5r41LedYt5ZztQ8jUl
nQiHQDCUBe9NeCquqqPRet2z+M+5PeX6fJtedAnB6zArjiS6vwRAKmaAHTSsKaRP
M0r+EIQQasKf1b/opPUw2aPGTvQHBSvM44/lQeuJV+64CO3Nlx/3CZNi3z35X3Wh
+Z+71w9lHFrKDIQ+VUreccXZNI4+tWNNM5WKjQKxOiUOj38Yo3+FANjPDB52cwEF
MK7LNiMUHAwrXwkSSAidB6Q+wn47nALamR1RgWg2jRRPbHhED33/BzTn+tinLnDQ
ugEBIwTMdhHMz2pEzdY5ub4TKpb+kWe5RRg35YEUw6PQ1ky2d4YGF5F4om5POYpw
9uPrJEu3Dhu2q6b/2Yt4F0TrxmSRd3woy7Kp5e7dUCGXWlNftBnpPfQdK+AWQJ1S
GJHohNCt6bvPo0ibXmKIMcciwMXYg/BotUhxfMxFuWD3APHC8XF6B79C11WL/WdB
xHLTp+qOdojj4sgKenw9S7pKCVjK+mH3LSwIYx1ShmD9OscTQ9XnOq59MsTMUCJE
ofwwg5P61PQKHX87XFhi0NVvNZludOfAfSqwpxWb3yR9s54WPTCXRFGkiabj186h
4KPoCN4ylonhfOTshQDivoQBIg0Wc9ENJW08chgLmkUNdRivirQ+EYcPzZTtqWDN
eVIFgryhe55+KOlry5ouvYdN3YPTzzjI2uOyZhvDGcymSOUG06mdU4IcHSaaWfd9
1fSAMFSPmNFyVUEYUPLyjPRotuNGm3bi7cq3VfNdWELzyY9S4t+IZG9l3x8q+Wfx
+l49kMUHtJobFnhmtKd86L8FJkr82XCUp4uGxDwoAok3jOUqkKMhmjuiYp6680nT
4bYMNhUAMrR9yeXXd3EQyALu/xLbA96LL8cHAbWslSyJQEhcwEzck43Ed30eq5Ne
`protect END_PROTECTED
