`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Osqv/20xDHpjDpqTeQYdEsVUca7gJo/+QsgQfa5WYbvZfSADWM5hen0RkiV0BqTS
KruKbmcckTGeUk9YBNOS3C8CqwED6wUHQ09bGUjx9h5w6MHruAOF41P2TWBMGtti
LTB8GDHQ4I5CLlBGyCq3ot9iTzPP5kkXgUmoVNP+pnXoSkV8Mii8MusN5aKwQUZw
ZfY8IDrHov4TZlXaFI6PZlkgfJE33gW7sAwspcWwU7PPFrS9tZ93o15AudtL5wCB
TUFbHA0lt+eXJyPKO3fphpc5/S9q/ppwqb7xulW2ZHgOkco1ryAo/+CHZxjXxGGY
LcFwrHlkeBq3Tnv88RAagXVFr4ViPsC2R2dwpZ+vLD6jHjGBDwnFgQf3pP+MAjY6
1ikPJc0TraUfaXFAWWrsvPVR7KrEPrDaJH3V3al6d727THmoPTXB2Kpb+k5dpUfH
+yYutUKBmbySvlEbSDtc0VWAvvRejNKHW5kArYExsv2ZZuWk3q9FMTy1bek1Dujp
NYJIUkqSnS+9JC7LQ8zSYUNyN1Mq8TOqMi9q5N9/NPyTxCqniQUFA8rn+0gxMguF
/g45aLXoCVSQwca8wfg/+MzXAeCJ3jmuvyWF6KGXD5jl09MUK9KSu3oe/gvSRZb6
PshhxqEHIXjjxIH5x9yKUOArzv87d4bUSqKXvEXX+G+YheAqlS/N4Y4EDEYaTjzW
KgSWJinhcgtyPow3ZsRtHsENCsDjS0kqTJKx8QMlpFb0lP1pTlPQnXasBrUgcVXN
uxbbWmQjAfVAqzwvHFWhawWkl0XUSSr4q8dsgt880H4Un1gFmVi79mqdhh1KuxJQ
HNhG4c3En/bv/4inQv9hKlK3x84811TmII4tqhODA8NAIRdBv5QTwnxcALuNfwBE
c6TyvV12sy+LK8OcAfVVftdsq7/pIy8EbQdSpn6aH1bzMmi72Go0N5YA00lKefjE
RQyKXHbO5RRivWjzRDJeEYczP9GvIYLPjUr760dAT/e9yOTUPmn5mpR/BQ+duucm
fUsdn6XWg5lJLv3ZO3I0V8r4Mip+33yQJD0orkDPrP32c06rkAfm8+EoDel2eFCf
Fzvd7m5PGyl+lhKUYhjYaedM7xRQtR+wIffXTTsbclOZ3ykGLIxSfXXh3RLtPn4f
SrtqZVjvky6MNX8ljPr6E4N5IQ8/8ekWmaFsTtHKETgfolTK9zhNtTLN2xzIfPsh
ufrjS3qs1kvgysT2OQfZ/4XGLgZHPw0HxoNL59aFyC9ApMTXEvZI1OiyBKJRsu9R
dfX9uf0AEdl6PtL97kNlYQng68TlqnKp8UzA38+oaGoxd21ziBIFocTwMZIZ+aAa
1+Q3p3/UHKtMgxfwVgvy8gIX2KXRYeAxcGNm4NIzKVE2EDarv3VEOuiiZLdBs5PG
dZZdXPxgzqgZ2pUpkhgv3MBUlnGhMlK3OAgl5c+rPQE2zsGi1jfOtqVoth8T9Hxc
1lPM7lZapKX9UYvjqjs7IG//kIxOKIUcUV09jloT1AQAAUBV4YBE7/17LKn+Neti
VpCToIjTbE7DosIuwNC7MpAXvP+U9GUGKhH6TNtQMVnkyTLzZRt4nJTyRspY0nkD
ru2xTPtw2fy+BmHh1+MUFMOi7rRi+vd8aTu38ganyNdT9/HiGMAvzjaywSDvXp+n
9LxcaKqLaSl+1GMkYOlsW4cYtZXxmjlAGPktD45PrUHRhNb+dL3t0J8ILFGDrGAs
gVMaZodQplnSu/IRpdqWJCMCyUFAta3Eqcalaa1+HpWBImgOzV/7SThgCwCZ1atS
vkXsz1DxOsoja051jKgxWisjyvd3oKJ3vIJsLcsEM2gpDqXgLYkkz9LsvZRmpgZj
UA214GHrC5RjOQZZHoDrkZQqXrXS6qXJIkct+HFSN8AlNnAdsBHFT5jIw3S2w8+4
IzOBIl8dyugVn9cIco8ENfTdHchU/8fFZW2O2CKGvQFlGaSL9FmZWBrbVRaMwILN
Buqd7YtBJNjccIQiawEAR5kWeC6NRTOjjjZVjZ0konPgzwnDtQ8C5isOyzAQzdEj
KJ3czmlJ1l1IDkChFLupucj6cHAVxFedbSNzyFAzT3iIYrDJJVbHkcGeUNBZ0KCX
8HCXQ0LIndzaqooBfvYsUJkKCO1gghRKrvJc6eVcvihpjL1keMlXsikySKIl/WSZ
bejofpza+6jjaJeA7MYKsO9cphM0R69yiQzoMAg8mVRefC4fkaqUXSRbHITpWraO
z68Rvfx4bYDAsZ3sy20hPBkmuCT+w1impuNGiW8XkDR5S4ixl7/N7lBqdhkAcxG+
Jm7BBZ+bUd2aW0sqKM/WrKMnQS1JLhyp8TLguAYj8D0BQNg4DuU0Y/Asz+19DiqN
TmaQCkjGHs+pcbIFz5NdFT5Wh0eoYiTvcIcZefu/Pdl5OwUrMQWwbXUZavTkS71w
Zkx6x1GvRB0HhzY80HQ4dkoHmPFek2D6ZTSUdDfFt+NO4+4hT+LLYLVWPgr0Yf1L
LnqWBpKLIZVNLgm1K7yuYehH8ipi30mXVd3ufae73S1VZ05lffuyklVpwXDTU2o5
odcAy2EqNmsH43Xz91oufawUQNnYqjEeQKZSKSBJt0RKkfCj8b5tO90kjorQ9MYC
QP/Lj1Auu2ea+VDkgZ1Ti28goPuR7E0JIjj/DprczPqJ/O/KciHotY4+484cXwzY
H5T6bZZAt0Fue9pmfnMWXPJ3pQN0CzZ24sY7q0RiR/u8EbHdUd4s3QwKA8rM+QOx
BKxuM+0BsT7sBWl6tEgGu09NrFYU772INVltfvU0AU8OaNs2hAt/HSnBraV1a/mA
7kiM2VTrQcg/zuegaIxLw4Zg0pnCauBwVUeB+O5yCUTuJvdeWmrVZ2Em4neUeAOP
f9Pfk/BCUf5YbhtLq8Y52Q3CQLGLgrxJphyj5wNRXjDGc4TI2ryhySa0vIlAfojZ
NAiKqqNA0UEWoWD4yQ4srLrAsepJSxK1jq1IQk4Gjt7PF08FROBhkfS0ogyST5f3
x354M11Y38JZ5E1uk10gLaCRl5933xWxdlRDHXVRokYiyA0ivhKCXS/L/yYiwoco
y557VF5OvIbbc8VRJ4i0aq8FwmfqWa97WuueZqPRUkLCEJfZLclS67UDs/m70Md8
wtpKvAO1SwwZvWFrJJuzvonX0seSM0iG90RIBo+1c8uDrcgdWTEyl5ZZlhDxw1RQ
zdBvW8gTz1mfVV9yihkqZJNzZFN2tC8xmUQO0UYMf8Afu3yzXBen7U7p8cKzCbMH
J/5ql8/bS+cVyqiVJc9m7l7lPRcuVAwPDEdNZ9MP3Z8jEuJDW6lRNGyYdGSvJyc+
vWzJ4FI8w1n/SyyW0XjzDc6yUUC8n4svA7hYxR6IkcQgqfaxGK8tdJVlKKh0inyN
0Fn7mFpsIx/Zw9vci4FBf6wprQDqk0qU+KY1wlIBtjtsmMZdgnUCfNER3ghlVNAc
9BnHx2JLWjH9y8hjt08xTTLjsHB+L52r9KxT79GK3FvNolWkZrpOAN1IdtJt8+a7
09M5UpWsQKLQIBfCjvKpVlyPsx0/rHNDzD+Zg64cxGOLU9ekKPazE2JYm8jU2Me1
+3WZ8OqYRIZyvAAtrYQE24Fvnl/tOGBMrgF/zlT21lpTVgvcmsZSs2dLFFlMEh+5
ReZ8wLlFPt+pGl5GgiSYOEkQKNJSpEwXjvlytMFBCnVQQOgVjuqmjKiJO793HQiP
EK+iPMHey9CFULpGuG+QnScFdtyhjVV/tiA/fvR8RSUOnVd3CU/95dCYvCAFwXt1
kkgbjZ71HYFtconeHlAvp00NmlZpGFHO42NxLcUn5Rk/c6M9QdQOA4zFLf1PUH76
nGD70clPgNnVkOyQwTXFw6+4QlYeieGTl6NtjiJgq/Uo4/UZXenFG7MsPkJ7z7s4
1rpnJAIboK7Mfe5jkHaNLAxv/Ti+38NW+a++zng3PmPGMy9qSWMMPqUTyfMmDyLX
CSAUoUDakp3gK6llRoY2OToNZcOBebWEeXmhitf7Tn2GT61xFbXRidg0g1N5jpmj
gZirOCVZc9Fvp6FJ0q83hjUeCERW7GiHjvtHuk3uGyKE7jtC41oVj7U2127kLVIj
P3UL10/5Fl0Pfr8SguY5AsuO1JI8ODsX2BsID982TbDvcWa/hwDICo7riWhlhsYJ
ByzV9kS2h2BD/NBdKDX1xLQjL9I7vlhM3LLE03yrSqcbc9b2Tv1ZIVGVdE8f39nI
nxoxPypNs5w9rY+vPGSvmfvZcWxHQlPhALkxpWq+EDqch+Jf5lz75XHCtgI9seRt
26mGKmtAWU+oHJhN/0/038J/eL/J7Lg+hI5Ioi1R8NH7wVpXL+Z/8xQukaw0IE/A
WZ+QNmh5aOKMhm3MremDCtFNBK7TnH+/z9aFPfFCoqWCFGaEh2Si52qeYMaqzITh
24Nh8rGezU9AAQXTM1Ido3Z7Qw/ytH1hWD868NGbiyP/5OEjHUoEQ1TnKP4aNokX
ITLpVqKPe+ynOYyxZijkX/15lR4+TMqpU9TQiRpyXF3kJ6ZkUZhdRO+40t4hHm/s
ZRx5xDgUgCi7FWgQ+PwwMQ09ltLgHNAGYQgtcxKV58fzMTQAE3qlUO7BuuUkd+5R
dq03JlOO15P0aQzOPHMcRGxahPCBPtJRozvjCLb9DHDOoobuxH8zIlgR3oWDPOg9
eCu4SudOhC8Bu6h+oDnNbta2AVPNA7YHhU42gVNQGOI1CChLRiSgHiMoS5IvfMJH
zqFvOYe0LQ6SzX07p5XBMMsefpHmn3twGtQrnkL8tAOAGlt5PITdzwdqyNzEKfA3
S0p4t3QhbhUcwtd+qT/0maQBiXPv7VBahA1/py9igs/jxs5rXfamX0MZJ3h/a4Kp
Y/O6o1jLyc8l2tCk6yq6GJ1PLRYWLUjOErW5ktUxeOvsWvtm0vNxAyTaZJE0RqN/
Ff6n1ep8ORm2Ebg7d2d50YlXqVdrQUoyEfsyZxhfS9Si14hkIU6wnj/1XXcSb0I2
p6eZFpO+IzMaj7/LLjiMrw3OHOfGxsy02SaBxyIn6ZA8RlBkRKyYsj1Vf7YjCdYw
SXsWmw1hwIFIBXmTq3Jz+xcc8Ea60SUJKNZ3gUXTsZSa56MRwstaermrF8LD+rft
G6ZhrQ1Mlsl61jBC2hx841oOpqOD4N7hEmvolcrQcai4faT42FWUha6xtpsmTCXz
ZFt84jXm+DVR+MMnfIqqiqxtkKjh2McVG7DkB0UVfgjINuwlPrfYOERxTBoYr5kn
jA79kaL+e1TDjxJAg8sJWnAXJhk7fqZPUCUJ0in0lfsStqlk+GTE0tB6lseVu8Yg
5n5kkEwlxE2twNHybCAF7p55sTIebIuuwTux0JLMzChfmd+KyUm7KVV6R6NlD1UK
/9kyDWs4jIuA004cfe+MiKYbLjN7S9vh+Yd6TKUO8Cza4LmstlJUzy4efkAA61F0
c2+UI98JfUYnm6BcnjWcb4M1WMszDeZKVvkTJuUVs9Gh5mO998i0yUrAKEMGVBGN
zraZQVTHOpklC0Cn2KEUOTcYdq+XYXdfeKm63/iXgymna9N+bxZfl8K3RNUH5Onx
qyjtb6Mst4doEHSEEhXsD0QrBrkswy0rT9fqgiR6up+fhG1w1Ksm8C5cRzDGBq51
HH+3tcfollNA50k5pMi31Xc40GWjT+xELMXWqlpuqvmDsY3j2Rk7q6HOX51yh8Kc
+FknqGDdqaBHoURa+h4ot4LY5+V2LYIJ8G4AUthKIVHuNhFlO1tVrIB0JtU1tOo8
dpTLq1MHIQuTnuFTb+50197Z5kw2ZODdV2D/4tSieJEQt/WqOthrhA6yObOIJ1/K
35e6TzrCLhpJNOrSDDVzbZ1rPW2at8J9I0NQmwkjM8wQ8Ec7bkxvQW3HVGxflgOo
FjI/IpbU6/BpiHMVpZUu3kBSv+ATwkJ4mx8y5e1sjQsSLm9ftXx4HSDpF/YmZBB4
759A+hv0RJtcn7lS9Z8Sj6L5mfBy+SkViNfRlbWHCwHH2gQQJydSiaoUQQTZtWfI
l7Djezmgfc79+kWOiPw6V2E2Yxa6aOeLE+HoX0QtMjFV1KpSmRFOKYA3X4EBhHQk
/pJFDA/HmXYMrFReS/2blM8c5KU8colmSQqL3rBIbNda/63JgzHojwtgUslGm3/g
5K65kJkxaSLVLqIoLso0iJikqQCxvA5w7ZHw5rIF7pZfUzCV9Foz2oecCKg/7Av1
6NE71eBI4bAkKp3plrURKQeC8X6wUDn1zhHN0d/btVXNst4NB5r2FStk3fuottOL
cdp+G9nwPFt3mkQXrd7PcolTVDaDmeBPOxVVucoto/wHQZNHoDjvWcjXTMjVwAMS
oRM5GLDZIv+GRR+CLPTVmpY6rvl/TX3qhA7/lrgNv6vEFeKc2BZ8/kAqbFItLDAC
cZ2t4AesaV03OpYxVnP41X4HO7gIoOecO48/QM2qb5E+0qfmrifhQbc52hUA/ZQM
QxqiQ+7ycTR8IcPtNvUlH2deJhkT+lO5iAvNblV+WLjXV7tP3SkYJ92EP+LYqDtI
8gumZxJMasjh+02nXObwpoa28cPvEOHCfyoWXyQ7J10oH4TwR9tHuxBeuozT1wBS
1LiG6a5FVAYcUuLWhzu5KL8WKNtQ4o0PzQWMg0Lk+5WvRc3OsJy54uYXW844fx+d
ucuF380Ri8JrIqNz+gyviTmXw5cGXo2kWml7vN7g/ls=
`protect END_PROTECTED
