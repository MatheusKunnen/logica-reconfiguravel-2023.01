`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NwN/G9es2uUe3gJw6pXyNG2Mov5IBa06kL3W/5nNRfk/+tzTARV9gaQqKl1iJ8ru
6hLmlZxRqGoqFs34qjO0D1a7oZOoJt0iBIvId0yMVn9L54Z91t3nbYZCNKs6ymOn
6jWzOcFjG6u8ytcaDHxbOv2CUKELe4QAbsqDvP5yb5t+ZVGhWHiEPE2FPpaOxxRn
GNIKd13Qn81TMkfvh3iziUdi9I9hNP6fcAtDeWOpIzfvecGqqStp5vtGBjHUGaBo
FTvT8yAuOqjBYroqc6I10ElhGYujZFwhqlS2sA8am12wnPG8BGMU3aSjqae3D9jO
12BK9xv5WCCqECSytqh3Pe4mk0I8m0ZqtHZcGoPIecMPtsBAgrJfhPZyIKNvGPhQ
nlwcjNYxKLT6O3hDf5HqC0ZqlRq7MhkpTpKuPL62kLCY1oD/NrXan8k+Dz9JpU04
XVX/pqGfwk38eEEAtyM60BxA4SQs+D1/IkxkmJ7wMBPYx/R05boQUFX+EofgsVgW
cAi/a5TvEA6nBLa/6C5J6rv5oFlHBOdyBJCiSn8mwqMUEFHpNhyvsDak1MU8zj/v
4qEUIwVETSdj0waIBL5lYV18BoEK7N81K5ZE2Kcyuo4enCMewAZprpW4kAU0T4v/
5Gk6LZnEA3HbKlGLoqT21uj2zi78FZ7lV0gSCJHftCdVIFik4Nu2WztqR/ZfBQO1
kh9YwingdRlMxUfce7Wxpu2dkZElBG8dNYXMjD4VuEodzqhvwkItdNDysPNrrRlL
/1Q37jc/fmGrguirKeiv9Oq0CGPZCc3ZuWaTz/iFD+YXzA/7HZ8ddQsFWDG74mtd
5VhM6i6Ff6N98kEshbipuAFcYGei/k6Txpa3pJdfPRZZpKX112ZKihTf+UlCDYM6
Dj9ZPpu4oiVv494WQ6H1VNJghTG+CaO5c7F3UVoWQLxIWz+kXTJTSF/iZzUyJA/X
Ebej04kRAAUwd5QE0DvPkADw/5yyLv7hMUfXs0rTd1sRQb5/ugwnKKFQ1DobP8rL
wbMyalB5Ra+Gd5zVPZZ7RT/c0CzEOgYtO2a9AnKNnGZoUDVVU8/Vjw2v2QQvOQme
DxPtfIlKHZEV6ksD94IMinlwsZLj+Y0jjFdjsx36Q1siisMgbnNtjNUgrEBM8/su
IUNYU+kI3Tw9IPNuN6vDKtH5kL1OOzCVTUqeVnG7UNGjthQ1HIb3KFjGFxXQTYKM
8wf0veBa4FWxT2dXiEHHWcwIqbrVaRNJtl1xaWJsQPDKeTo+NpQAHvcLIktXzTNi
n++fva6Xv6tysoii9IZymBLwjaBtqlm059y643PxemxzRxrk3yuOuU6EDBC7kC7d
sCDpicJvqEQHhLGHDPrFbUrLj2kbV5uuZV7rhzVFAIBL4Xo6FOsJOwvzj9PCLon3
snvTrrY+ywdGQ+YBg+7VX0PuAqLgqUn/ijSwlQrp/joc+a19y3PgEy1qpxVxSjMf
i82ucQj3V3omldaCh8/joGjrGoNiP0797v7WZhfGZMAYQLd+bOL32pL4GDay9AtE
kEcfk0XxBd4IAKQsF9QJvLU4enn7urkOJL7G8Y9Ddvat9NCjVP2IbEr7oCrJM0pj
BvUs4lEcPgmZB3UNXS+x/RPhFvbc0YmFt1zOkeYzFyTgly9GSzB4pf2B4wD9UrrB
TK3mWrHV2tRvFktpqIEvp9DnEmCYc5f1m4C0zUWU1QQtgx2sh4T0fJEPBnybt5Io
8Tk/6ARkqcb9fBvafA7nTAz2ei+pD1FaZmeTVoSFgPUwewLQemu7grfdH8Lt81MH
VA8GFtsf2ydmutrHxQmg8Wa3R3//+ubjTy7yVP8c2/hBsbslrxDdj9xCpCpGGGvt
EUGeG/XPaqxAwvescdymJvFVi7DwjT8x5xJsG71+C6LPLz8OR4PSe8oAqFQpcfsh
9716qeBRVU91/uBs5TrUzIc47aW0LkfBK7WP8QNyd5K0OTyZw74E9YCZ9I1UaeGC
jetzZEqatxpZ0o8MrkCKdw==
`protect END_PROTECTED
