`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mnPqZAnb2BfhJ7yLtxASBE2LJadl74c5f3fjzBshTmA48yTXJkyke0q9TGINbBhz
T+vHi5wjeqQoZZSVJe0TPDrdHLRdqIb+r0uDjSHKbEEvXDMCDJ3AhbYPLUmSmNeE
vNgvL7NgS7y4CUo9mh+mdmXGF+Z7a+JVm5J2zC6YD5N9b1oJvsRiiCANTRZXFXPf
+m+GsTXTC+FwQUj+K3UBA7ps/HEtYESxvPijhwuXMiT3pP7/7FAbtS/vJAh/+RnX
KduhaV1hQV+nlDZZ5c06X/Gl1w58r3UUPxinMIkMZw9vVniAbXH/MqaDDsvAKhqt
orYYwpe1p65LT1KB7szYCKTtCA6tJR/a26JBVKdPGYwKsZkguLRdab1+bfreucqn
g2I/aO0LPZCuSK5iHbJmR4z4NAtDo3uCq8s1ILjfjPWtjRjyFotPnTODvGwrr0f4
W3GszIYME/i+BUxZJ6IgDa2aKrst2g5FNUEOE6q5QGzfRpBZZLIFnxDpz7+/7FGg
5NjViXYtmhAZB/SpxIUHHXka76fbNSyZLcJFq2WA4gRAjQgEEjg4LuJG4XJlJGj2
QXeWuG1AlyWjluH4lXyK/1W9nUdnYahFe9/5cTRNdCOy6Qkjbwqk3qV0LxHvP+4j
KXGMyomq2PqXee4zEOQtFSwDX6QkUJ7IeBSohjHrEtzNHr50Makdhpi9EBY5bZZB
Zd2WVaI4vp5bbMa0c9i3uL7wbUmZOVR7FpjuoanKnv4nWvGxnC29zW7EO/qCtuH+
i9Ph8MDCXNjyq0jYUKQXsx5M2aVuz71MjwjpBl085Eb51c1HVG9x1Dh4XkcfyeOm
li0q3nBUFisK/ZZG8xRxaIHZjL7iO9lyfndC9T90zzS92hFYjghlUISbdKn2wSsO
33LFVrgW3mtd2ltfkxqb1tE043zJgupia6LnM5pQ35bzUa6ay/2fWVP8W65rJUNe
+mq6RVP5pmhNtBEFY71FH6S1+hfXxngtSnWlI6B3FVF2h6NfU8RsscX87D+s90tI
2IC9DRdoMD9qbzNhazqexQUz3OfBIef88u9X4iSc/wpdrHH3AtYYcuiv5YQwQzsb
4OfvZl0hqZHNO2syaIT47bY0edtiU2ZBvni3mkeEyHSyxlSBd5SOsDcSKolekFgd
p0f6C/CbBBWEv048U3XSYTC8EYqMHIhoJHTCDYFNvXj150quKqlM3O0Dkm24+mzY
7A0UzOWx+1LNCxcGhxEe1+mXn3nLC2kB0LxULlb/5f10ItB3XIq8kVSSm7BPVG8n
KH5pZyJHuLzCopqWuFRmQn88yb9GVSyKHRf+67lsfI4btViG9GLJVtiwwRFSLN1m
EuM251XpWiSiFvyvd1Gs+ENkAFgFaA5Sn8iBHaG/iFVG/rcMz4YAIf3z23JBEZSR
IwNWDCy+mcpJz8l6X7DQi2buppO5LwC1mJ1kBEEWSA2pkxozbWimToPlv7sZmuas
tX2+jRs8sr+Mv2IYkySJ2QPYJYUACp70Jqcd9nNy3VzrHioCzvpV768gvQDBQ1Cq
gH3AySchOOyQLbxJY2jSXu0aErkfPJspf5xAwCsV2Tx/Te/JKXNbn9syE41cBM59
GsehUzbx7rOT+QbQFEGqHY/dKoz6WXAeY7IH/D+vzRQR1tvRFgGDHwuLDusIS36S
3c04yU/RBEL2Ime3yiUQYqghXXuvm4xtYCHCeMCfoDr2Ul807PLmE+WNGXe4CvmG
H1CWcLDCROGhLLVPEmd7ntq3RnrdSVGFx5vQ1PBR1kZk6riR3PqTkCh872rrfHUA
txkDmCsrwMlKtOe83uwD54xU/1PZLw5AU9dQqd4uSBJ8lljnUKYfAmrLQ4G8/k+D
cjYqUpZU1iRSo8EewdMYvwlRU0K4jx6oZx+mzbGudrH/Ckfwkl5o58Zn+jMAgdIy
b+ooPDNzC7TP34PJVmveUlraRLSPw7uFuNXaRxG2occx+f6BqcAFbPCvuohrjIYe
thgDuBR+auFOad6z8y4LeY9zeE0SJOcLSDyEe2E/LH4JNpE9BxzInSVgSI3X0o23
I0DOHYCr2uungKPg3V7khbasK99EhGsIgrqD+1AtRbnfn5MydnVkzZBCU8gPGbsn
QpBKtqLoiscBQm7tfbkOVwDzmxUPLVTvk+dHgj6bLHRKeTna/0PXmw39RVtJfRF0
PCpHnPCNevb1zuYIoMBY4PFfxjI/3OvaDzqoRBNk9mrSlemocEEWKAaSkZmL0iZg
0UD2QIHp1+vdBub/s5qwggNdQxLJZieMUHsBQ2BfyQZWPhnJOKyLy8tDKORxAfF2
dLKbzp2x+ylGjk8YEI2+gWcva0Y/vifPRuFPIvGi6xar1XUYlmS/epv6rthqzxxj
2qEZHe4sa/ZA8tD5UZzdd07I6HTsTpcVqMQYroYm06PbIK4tlNC3+R84nlxw/w7k
NJ8tv9hrVXl4YfOwQ1p3tjSxF0uRpwKDaNdEabFVgIPJ3N2TUHnCB+LUW+x5pTh/
D0hrC0eq2IByd0tn5kfKm8rz/8KaNL9dVjZDGR5nJgUMYVfSBikk67EnKlPtnmiG
7SWbE1Men7b4EPF0I+c1jN/gyaklwQgksVjEJhOmh24z/0vqd7Rfl+LTqmpgbUT4
6C07/7cdbL2CvlNHinfEvBBnp7RCLu7E9R+ek/Q5pnR7K//LTaTnsjPM5BphQzrB
5ZcXSoQFkWWM53PW5fgOt8Wjzwt+E61wCQlX/03BoDJFQqEuyv010SprJHlWqfQZ
K/+DsyoKVzS7OjhDr9ZPoXfARn9dlz3tyup2Ax2BOsbWuwTB0rjUxoYzAnjK0Gc9
1hT1JOUVo0SkLpgsoVzhLIg+8n3UIU+CO+BKDgf99KyXeLkgiKLtpQDZREhLuBQy
ADg8lhT+w8fimRmkH+JH8SXj+YxeBRqxsp1drcRbzcBYv/QSXTMUNdF5Ogn73AzJ
ZvVr8ael15vE+y01Tk++fn+eYpv1nw/FdBnCIzGYMUAzk6PEW3KQzK5Mlv0x94AH
he6Q792VzY4+AIx8gNxLg9uqVDYFmd479icWjNH2TJsvF+AB4s7jD+VBwkaBu1Bm
Qik6/Bx4gMi945qOBk4U4cSAlVComkFRV8m1FVrNj5tgjpSxYEHsH2gl6m57Hp8O
SNfJ0NO3uSo+NQ1IIJ3U28EOX04lzpIBdSbNwR0MNg7y3XNkFQIe85pZwemQc/j6
lKl7yh5f0UlbqVmHVu2Wnc1aOfsHg+ko/3mzIz9gA9WUbjdfXajm/fB1ENiCQfFZ
5bcFVteVy+iZLo1Hshbc4wx+GroULAh6tbjizDo7cgGX4rO3W9Dt/0ebbpXeEEdA
bohNIdcwPfTxD1QZH7JcO0pN9g0ggpwXgktJ1Y1+bZ0QngsRcVGns/zCvhredxVg
i/DDJW0MDWV1NjKTSYVv8xpvYQ8LGJDrYp5vIEy5VYA8fQx1I5TfTvK++MUat0Je
YzgdJRIIH9iF0F1MkSgPR423Cv6gC0nTVCIgHVUE+3dxOdnpLna3c+lZcKiIyoks
i/j3cVFzyYhybqiL9Q3CWHUwcy2OzO3kwlkqsYDH4kcoJtJAV0x1lirKPyLLdMZ9
lT1vNu34Xvj42c2VKp1uP1/qIzYj0BzS6YZACoCaZ4D+LTy3BrYKsTY57B1A8dvq
SkFDd9Y2FCgJgvwM1Q7xYuxVduWUK2MLDmZfWFLxzltzILNMdtLwYyy5rsM33u+Z
1FtWm/ocwple2BOO0wpXeKr4HE9nBfVsxpENyc5tXsm6otQscOGTRmH00XS3sSSf
IUfvQ6lATSJXJx8wT3eIO1CkWtNVlIC8udPkfc0w0yyVQkKq1SSKnfYSacIUN/j/
DAoJrqbnJvrFr7swSG7pVc9nC7zexvdpcPcXJzFfQBooXKuvzZn3bzqP83C4D9Ho
M/6PeZAwd+PjOzrvKzpevR7obCGHEn0qnLm0qcK5cVw9GrK87wNlmTbbi1HKkcYI
NdE+PIyjkQnveD8RnkkaAfoDq+eRcqwDe3i28Io0ryH/LwUpLEuRi4eey9lyqMl4
9pSp+Hd1qkn6DkTt0nuYgOo0PHpKJxUfJktg0xa0xF/k0hTMUfSzMqkLbAhlqBTC
OoIcLjsxr8vye/SIJ4Ky7dfBKfdIhfKeZ+MdBq4VVIEi3KbnykNQDXL7/qEA1qAh
NgF6KESDpS94D4AYsCGGU8JDr+gZHgEbRtHgrNTTRKBpwODdhfKJPkZ2TLKPO5dc
qHyziZbA3/OlV4DLsgQXNz0XX58QMHUnU+rq6dpWkGvhUIlGMrC5dOAOSZJ9jIxg
yAjK6qUJ84Tw4AI3MNc0hhiK4bK/HJfYIX2FjzSNkCG3Inzhu5337q7yEceS+5XQ
GwwK4XR+ahF+5O3G4Omb+MAZjyrz/bkkWZ7OcpDmzaV+EFxU6555trZOdM/0hXD1
YbsaVnd0CopBt6oIKAXP5N0bSFlYXfxPr3JiQFwdq0B+hr52ysolD32BBOyoXill
Zv7qLTtntQlEhWyDGR4MnGEDyhckL+hZKZ6soabvkGOYSVcpSpXuublQ5z+0aVjS
/qM2K2gbOcJQnQV8WUYJo5ABM1m5xzHStwK+7wAI1IU15sZejS+f6Ls126QQnx47
UUQAW1I9cRBhtzUHVlrplIPfM0EFvrKziUKXvWXRpo4LfQ+HG10BLlXVow1N6/OL
QgQtEp/qqiUp74rKVc/XiyhnjBmOPEIn0dccHmbyG6aUemiyQb1wPNyrBaV/cVIW
WXxSa3GwbFeYe7XLvzAveJJ/1f/Gt/9eCDqtTcAuqmxJh4wVeBqSGBxVjdXz4iVP
loydsQ6IIbQm71EmegYsPmcrNtfFpal3gXTrFdaUCJOfkzCPHnaIJIZVy8mWbjAf
xijM1NMB73uJSRcodbmbiHglua5z6T0VQ6zcZwP+CDmqEFW8rzbl7XMh2IGHsQTe
AWT9aOVcXOtKSTswgZfX2QpxfWljZiKMTdWqQIa4G7l+n/6Nhp7SOTgDxRCIVDQ6
JJvIdSb5sqfsTab0pEOiOvSeCdU5/yDS0jyjzJ0IdN+XyfAm8gvt3/IGV//Eo2CQ
HuLFWpOUVYNz3IrvoVTBFAQjActm5zey9F70y4bHRPJMjG207M3yWzYK+qtDG7Uu
WvXQKRFMNRqjpDdXZzKz8je7L+L8tT9pYa/fIaOPUqDPQZz/PlbW68GcgP2tF/T4
vzFodMT2tLFewgBEAZQDpiUCMuOLKZol9T+oEBgYzpGtmhD/EfqneyTIlwxO6NUe
1TOxapFd/G5CnA1dezPILenWumA4dyNKwDPsQyBYrNyr1IRblgOFEq+S+a7PeHmP
KhU+ZvLuNgkgAmfFukhWFIhxVhOB5CyGzsAsd6y6av1AqwpT94e59gY8fZvmlATt
rhMpuThunL6Boxv4Opa2zZCy4UwVkeiiGl+hfr48P6pt4Lrramb1siLNf/yXWuSk
q74WLLvAnyIEnJ8gfKkuzla+xlMe/LDKJ3ZYjVVnho3SAzkYZ+75ZQBy+69ujEOq
y6SoAH1pMX0Baofl0rIdjiuRKNCwQ5hO/cSiX7l3aNGwpog/mSqTwY0Mqa1GSzVC
GYwB3+sfVLPUh3crUTkX4a9I4vbIJhjDCqPiuVMaRux1+wHbkrvvPglm37P+3hS/
6uSQdqcxl5WhgZD+vmAUa56SdsT6o4Id0ZYEO16eIicvzUz9GLuBk+9MjjVpYI+B
hp3wsEz/IqWZKFbIiE6IwjrZl3NxTK/fqEJ+T/+JF32eueUZfLff6G9zxni81wFe
GvJlt3Rvpqg4cVy53lcHSsDOaWlUUImNCSKZ79yR7z6QjTil2ShrEczGwVncN5v8
g5icKKtkAFzHJc/sg18UwtJvTEPx02Ur6uc0k7FpuuCR+pYoQBCtjpKvhlsHvFE9
fvkn2A2B3d9GjuU+0vyCVmdVkyD3btfUghDjLUFKL0M3yyGEnctsUIS6CiYO0quU
4+s/+YFo2gcxb9TBpDnihntxInhY0cOQtDZF8wfrolqx8IbllgG2Hb+Dz4HvxNbl
fPRgWdrBagbwdiOSifus+xRf/SMIu9oV8PXuqrJvqrQ3QK8Uwv/lLrXLGGDSZ/UT
T+k8yyMwy+j5THAf+S4s7XWSGR1/7EMMCDSediHPCy9L9/3sna49CXVOn8gpA9lL
V2+C8eEVnAAgDMiPfrj8LRfhujVOBLSTDslunOxNhyxx6xX6DIAgEKtAD//mbaXV
1YCu9XrpFGhFppaCYIHpWOKp2KjTKq2g6kNX+0nSLvigejVv/XzwZfaS1G1fOJvY
G+f7nQuxyVm5LQPrbu/DCX18p/CwIzANAsSzAStX2ogdRhLHmwteCJKKL9uJDUOE
zpP3OGDUKBJgrtJUK5mFzw4pOlrmUvaR705UVpEBrmP+MLw3p6Joxf/c9V8E8jP1
IiFzKz5KVG8TyHlxkPdG398SmQrIs4zhCEswqNzrPty42yQvH2MpNauP1y36UD3u
E0nxzKEFu1iDpsc9npVQiSHfk0oDovYpTgjI3LiUzmGjTaNXaVb/8+Uik9wc44e1
eLleFzHpdtwhL9mMUcoOmTAEeCkgJCWzvh/lalxUfRTovoNQQKSmkUbo9oqlAWvv
eYy4DzUkTCxnyjFuZ8N2ffwX0XnW1HrOWZWP767vzCMQYlufM/Pbl5bPCPiJKKfV
ZnIveYzKTK0IezUEIk9LbLRBBlhviXxOouvskevpzXAEHGsBQOtuCr3DUxN1STju
v1pK5ZbskCc8R5d66yajmwcGTjybnrf8YbKqiOxW6CWGX4/EnlvQSpKwWVD5uVUB
lKMULDZtdeG28eSgTUfr9Vd/K3f236iww04JiKplKLucCi5qINDlZYYbP3xriov6
VfQVjx1lujUQSWWinO6HGON39REK46zb5AU//wZlL2BFHMeTFO7e4fO8KtZ3YmtQ
esyRrupsYn1LPgqVqtrmxEuiF2Th5q/OEcR2JcellcVYmwgDOFXaNPArgWQ+EUDv
43F5ufVpmISGVt05S91uzzGHQCYTAqkdTKaaKkBCDbOrYRm0aoR51C2UOyDpGA0K
FNGFDtYNNySuzusW3OCBAGx2HX0K6xMYQCqnNfdFRAE0lzVeqHQ6Eax1d1VZjTA4
wF72GOQsO5cdt/8DOtfKStPkzBSQF1O5cfP3e4qhs3djt/gm7FEzswS4jMPCcBe6
Pzf1WRPi5oPO0XTiXmTPI9TS6W9rY3wvfplt0jzar4lpnrPYBPI2vcCc28e91wjV
FL+y7VBPmhgbR8OdKNzlleojs1cYWzqCvGgDcnjCozHAmGD3j1/xRIS9a7D4qwjU
e2+QZgu5aK++pIyUA0Ix8yCVaYzzxDo2QtUP7tJ3fJTHtpay3mhpDF/h+9jqotNP
w8oKXb4rODRQ8LI/8G4lsTlW3LUWMs4oT35Anz/YPsNoQLVlPCA8PKOrdsMduFzI
sh8rtxhKlD+S6Ze4mncDaCvDvuNjbE6eEJRDy/P8BAgQznIuUjh1BYRrEd5c2z38
CD3DOx7uzBUND9eWmpushkkJkHkKlKK4wsAujoCt0HhNG8mmc145Psb30mr/Ixt3
Ne7vYMDGba888YFG2c7gldx20ugnp1DQoi2KuN5+YEMi9r+zhlcaHrf1PjnFCFxq
xrEL5HEYfNgBkDBDdRo4XwQ/FEzXV68t9rbTNdsPKpBFsafLp35TI7V4AIedkC0e
`protect END_PROTECTED
