`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+/xhHp6K7lA+TElf5iIwQh4xewmDlLT0A9CufMJqU58UPIh9vrx+0Z4wm76Q/haA
RthQ+FW3fKMbqqnNTtIa6xzYNJ8n/Rx+m23ninjdwdGa1qZmhhGoBWIbe8FdEnlQ
6RwyxEAG5k70kR/fNaeEpOAIseb0ImN23ciMQs7XUpElX31P+ic+B+14DX5SwxnP
EdnpRGJU2/adq8yKGMcc0sahl+DTt7kK7qt+JLz1GdKRMmCh42ia3hExs1vj8V1a
rFtvb9QadZrNYT3s9AVRW4u+7q2N3+o9Fr2TSlvQlwfpKIJ93eU+LudR6zU0Tv9o
1b3xQfst1fDrdcDfyGTKOVVXk/mds87BFI/bHi71y9/xEI11ZY6U59lRl8KP3Sl8
5P2RbHmgALGtbh3QG9yJfRFFhl9Jw1SGQfgNHI6kzty3M9i9G9+vZRzy0G7vXoYU
8TNWGABwW0CIkqxiOkajSJdcVd4sfAE6Bnt8awbBeQ0fg55QXF2Em4w9ZS9RYbrP
fCulg7R03ZDXwXlYLR+fJeBN2Y2Wb+fjgdk4ROpaSiOmvRcyZ18HXbBIICCyDNFl
0pIZtUP0hID1vuZIVWP9r1+WraXi4ahPb3tgPu2H3FJWk0DoJiJRsYPnRmWtEt3V
IELmnZzCgfnboVR80cXMHeuLuoDeFPwtj6oqK4B0E5T7L3+VjRMMnKgsZyjcR71m
V1oE0hOvphIfhXQGd9WunjJA3Q5kvO8aHhlkADvfnZs=
`protect END_PROTECTED
