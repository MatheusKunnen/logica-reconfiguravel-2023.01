`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B0Rv6dvmS8yS8Db5PdX8uj2JwRAqnE64ZXwxAKYfCMECBoj4O0qZE8q7hVBKayGl
ICvi7fq2S1jNKZmlxKI1lFTkU52vUReBH8rKk5NIWUV4RKdoROXwS1OwU6yxFstI
oa0W9vuIeeC8UCQKgz7kgeL9xOJj6R+APgpvwwH4BtKpKSD7m1HA3MjFEojDMmJ5
1/zP3+PHeYkMlpxARS4UcgRCpaICdOh1lXM+3iv20KPpsPKe5ifO8ktCVJgByit+
tzh6tahDqyC0hXiBsjt8RhGQ5RMYM3LwBjA+qripLoPZL2cU242iCZYdYs00mPTW
pAgLSKFU9T/lcLLR3dUDS8wZ4rC01qHqrmS6ojAvYOqjuty4jdc6a6iKsQQhkpkc
Kzn2ifz/u8K3wtn6K+RxYgCgKD0mlIX1/z+yV6X2WWtzSPx1wEk38qa3qd2Gf9zK
DTQW8pIG5XnfaLo/vDl8WSwU4m3WRQp0vneglPyKJXrEW3FgmqRiXuqcI/Pew4Zf
asWmOhbIpbg7Ky8Au1GVQUDq83u2TJzeoHOZYrgA8a6XBTRQ0mu+DxSV45yL0gpI
fLCVuoFcjpJd3Q7VxyQK5w2PVRjCNhOIkSmPdhxe1WTh6U9SdhsoYLuFJtoEykDd
QDpE5qyF6kCY+0zI1g/J6TFWTLLeDSJxC6FQT9GwfFrv5PuFtvl4l+q7fShucxfw
`protect END_PROTECTED
