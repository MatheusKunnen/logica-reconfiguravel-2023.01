`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M8Zfn4KMwPDsTemi959n/JtSss72SNXCDmbF2k4LP7jaW1xdXLgUfaYsqRhJJSLc
iSd5FZ3WUeUTbsWBr36tns69C/4KVrg5tz3Trw2qTcn7rsPZHXeTUl0cALcxweTP
lGB0m21ZlILgoXhTurvjrpMgyOGEDkGqhXxfmPulapKjV1poFejn2m9cT0HBDOnd
MbDGEOzGRCYpp30ivvIvVRp2rsNWadYsht9+ohbEfiBsGB79XLkNLn606IPaczYS
sBqDz0B9wGyUR4PtEkeMWL+xZiIY4aDlpTY38rELp4Nmm9fuqqVLFPvU+6alnGKC
wZlI73jhUETiN0GvmtWep3AepQyVL5NaVI/fF1p5r3NxqParK4bNtpu3nz179v5F
y247bF/YxySsfYbFdE12uWwPf0HCxVBXibQaM9yWQZjznoU0ADJJetAp30S34esY
zi7VP8zksNqO/Ylcecs0jBRhGE6ue0+wempJJQ6z42q5lCzqCn5fHy85AqvU571f
LUCDdhfcIMfY0wff4im7yzVJO6CUGnmAX1CfwUUgiCxX7yIPP9QZ4qko7HlTzZ8S
N5Z8QhVES30O4h3u9+ZB8OK4PH793SiiR6zBxb1IAbaIA/r25fZoj0DVZk6funi6
0mS5/3owhg/SM5KAGp/q8tzRMGobF7d5yjaBLcCwqR68Is3d25jx8VLvkuTMiXv1
TPNDbef0A89NMStBQVAW0C59MsWvd+0PHM0a8NZZHcBNkw/lVdwJ40AcBpvAgwBM
3EVM+nTE3flt/yWy3oE6VkbgjCjozZT649MrSfSsPP7f3gMCGBbjm4vljtdhjyb2
vg4LeSe1hyRqGbqRz3yFy2EqwHRlk2RQJiliGeoXftfLs2rfoWjW0IVByKNyiBDG
JYcF0ss1pWvHaPv4eBylF6tIJ0HGsn5g+pTkuhY3/MQ57QtxejgiUe4CaARptlTi
e3DDcdPzQAzA+gCXud6boRIG2dxlH2D3G9LOPVbiwX+7lU+HQF+kPUbPxjujiDnC
Cb3VkxpmvzXz9fs1xhSPokYsOC1hzYkGjJD41FnR5SjFp/Ucg0GwrTd1N1/4A3Ik
dIU++GK5jCIVJt5fyKRMtCkzS+dErCameGggKeicLQxUoBDvA7ZJBuyXB3U1ETDs
JFID2CB4hve5u5ktGxyxDa9DhWeqgdSobkuLARjgp/TR/rBwsJUWXSYnYIfMYs8/
hig/AAtsRuxIK7vlxd/feEmvJBHDGxkGgDgZ+mMmyqZJIT6OwGJB+N82UM0tfyPm
fvFvrqwGbU3Qq5vxslPrKHgcirkEhhTZwRYducNFdXXP35YQObAsm1QLhLLIaZsm
r1jXhq2+M+J2njrGQ3/hgbsP6LhX8CYByChIbERt0Mz7mLYcRKjsCpUKzwX7YNXp
gFrj7pL5c5NgNoiJhb017JFtmByXapYKvB24AqzQgq+DNUVJLd94xuFO/aA7OY0h
GYUqBkhvpb4coxMUh1LPIDDfRVIWKo2IFbMky6d07yWRLfNPWfkBkipDv7CfbsIG
825zYCiPJeJfj5V/6+0rFk310mzmDVEZa6fotDn6CxnRVEBqT0ZEkUgsjRd8K/gx
6BnOp4InbpA85XuFgHKGOklf7N/HgaOiG+VOlyp5vLEgnaMReyEPx5XFtbBCi/lE
D3ir/s5MkPUuktm35Fg6fpr9K8iO+rdny2j8FcP3ScI85fzNgVuCALPT0L9z0BPe
WgYNASr3U6gNJs/gFZaz+EQKC0vCcTWBgtrvny4RXCIAI+p2R7cbf/Aiw0mS7aPl
sjknuh+BqRHISYkPXd6C8pMrktCkD0OAvnz63JsOb3KeH5uaG2+g6nLYKd3h1C8I
ktMPMDdbXh5axU+xkjPDu6ZABiteQ9CCcPcY4PdDS6bQrQdKlS//f42UhROpfrK1
Vu0Vq4+CEdKfdeX96LQ+9xFPBxOWdSU+hovJxm2mjUnEEJxXslenpvQRmEP0u8Td
FGs9p6Jq6sAGB9n9E1vF0CXfQIDrTtU/WmyJVlw+EiVuquMaO/L9W3+pO5H2e1cg
DmVTL2u/e7nZ4qIuN9ZpBw==
`protect END_PROTECTED
