`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WA/rfOJeMOsyhnkBXS64dNIe5jpXSu/Pf4NXwT8OjHeCDoqIMnOy+mtZ44jjDh/A
3MtywlQXDeoVaHmKUHwRSN3QUIiHiqOaCDLH0WXkP3XFyn/XEOxARjLM8KgEdvsi
DzP9T1JxDcPXFg/+3nkIWuXz4DxnGVBz8FOdLHjTKEOdtjiPLOW2dAFAWiwtRPkT
Jz4ccz4Fsdj1RmBpuKJLPYozpQRQvGMHxGa9CKa/ZCXLBP6gsehWV2wCdyBIhcZV
DNWXP7HiY/qEQoUxA1v+RafE+sy/UZ/PCpjKk60rSUkPJMJznMh4sOQIcHQgmK0q
VlfZ8Amo6+Zu+mAmMlSQNcF7VQ0jD9uUnYfNBHEWDbZFSOGo5oX8U7IbRnTK3y8s
0N4jrQPl+ZbUPjzZUzlVd4r6S2g7E5UkcbSZJFYFSmKG+kruMrsVNp6oyJhVya3V
sswZ03fBneujAwWqvRpPLQxYYm77SYGpi6yt27XH/yy6ftq6dyubIh6CZKsTfAlH
btGh024dWe7UOLJGNGVSGOsExfbrbEhEtpzGw3/UBkl/B8HovdscLk9sbEMjn3Af
Pz5cyIC1+8bq69HEN0rdpOItkloGbZzKzD6eK+DX/Db8FH9VD/3wbw1+JfYOmXWi
kdMIpNz779yodJuF3ROVjoYJDYxgvM3l5X71FNE1/h6xwfxk5bTxJYT1chsP6/OA
17aLJ0tGJwHTYetaPc03bG7nP+oxCFapDD3ONK6UZmAb9zBLRtB5ePO/Vb778VwV
zLtDr6AsSs86e3IQU2sIkpIApLWX7bFdUhoNl+/pX6F3luejT6h8ZFt+QBqcf9yF
GHIv8+H8nNFAgIFW4gB1I9UO1sULqmRbt8M6PCVmf8Y0HNbGprKLAOe/CrCIpqbs
oNgnJKSs24MFiYsnfSIwZbei+B38LoHNlVPvGvpsOi+AFHPVbXoDwhabmyTum+ZT
rrCVHS3auHZjBTBpCoVKsgEEiY1/kUq6ker/o1A3LI+q8B6CEBMUSB1Nff2roJ9b
iTaRj1G9fAjOb1DOuPC/rf8LGjNLdzlnPDZ+hfsP3IT6gCPRTGJ0DiEh9aHb0U8k
qwZ+xtUMKyVjb8JDMDKp1myR8VnXz9GNvl9ZiXWoU0CSA5inRWiJG8M28eqMNkOI
M6I8wS0r8Uooglnmxn7s9uqAWqHeDH88Xn0EUKLsLc1q/w0W1hJPOFM4sDbUtBgP
wjtqXFpZ4wGV7c+qy1ymHDpiBg05Q9Ep3+0xphcBI/8=
`protect END_PROTECTED
