-- HostSystem_tb.vhd

-- Generated using ACDS version 13.0sp1 232 at 2023.05.10.22:16:57

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity HostSystem_tb is
end entity HostSystem_tb;

architecture rtl of HostSystem_tb is
	component HostSystem is
		port (
			reset_reset_n : in std_logic := 'X'; -- reset_n
			clk_clk       : in std_logic := 'X'  -- clk
		);
	end component HostSystem;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal hostsystem_inst_clk_bfm_clk_clk       : std_logic; -- HostSystem_inst_clk_bfm:clk -> [HostSystem_inst:clk_clk, HostSystem_inst_reset_bfm:clk]
	signal hostsystem_inst_reset_bfm_reset_reset : std_logic; -- HostSystem_inst_reset_bfm:reset -> HostSystem_inst:reset_reset_n

begin

	hostsystem_inst : component HostSystem
		port map (
			reset_reset_n => hostsystem_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk_clk       => hostsystem_inst_clk_bfm_clk_clk        --   clk.clk
		);

	hostsystem_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 25000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => hostsystem_inst_clk_bfm_clk_clk  -- clk.clk
		);

	hostsystem_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => hostsystem_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => hostsystem_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of HostSystem_tb
