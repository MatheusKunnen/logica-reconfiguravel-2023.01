`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1DB+346C2GrCDLKW7qdiLgkR8PKHZW6wb92lAzaxWD8OMqLweNo2Lk392B0JQC3n
HcEDbFFbwQq4DsQftGPucELpDf9I3e/9W1tiRni+EADOMcftHsCKFqrrjubxliWv
ewvTOy0zyKMVw1kgWVOO/N8+LtVksdwUTnPqXhj6uN4vcK+uGz6MXebz0rFkcyC+
8yGIEdcchl7wbjILjHHGGbRscs0rM6RDNdWWFDuqdOg2snujsYuplEah7nr+qqCQ
ZdSqKLfrcU8BzfCakIB3vWcTbVHC47lRsBnThCmlMUgma1Pk8fj4AfAFL2skrb3S
KmjSy7q2oR2DwhXaE2drm5FLd7MY2Vw48fM5cUFaaeRmBkH+WBNmG+YnrO1UdFYS
8FA8gpQYC8ueReNDRgfCcsy/O1ACrScE7AmOh362jzGGpfDfpD4h9/n0EMj78oM6
MP+R0TS2gq0q4fXiKnQ99IX1iIqpLvGuksc1VVsN2MKmz5MNKdphpvzarSIg6WuR
3Vv7T3cPDkaxUtFFDZEB6ZYwbq4G/e8o996YOB0EWQijUC+6UgL1Rn7CtuH6YqS9
okez84i/FDbxhEJuPKS2Q7ZzcdlE4ciKQlB358OvQ+ZB93GaruX5iEUxs+a277Sr
d6txWPwehM17FnJ6xo5cpqa2MeImJTITAEIkJh/HR8H7QCcLvkMkyjdCGWBvQ6DJ
kSy6cv3ZBeNEydwChvKBXobwrX8Dk9r7/OP1VWaPgmppBAItMBS2idxG5nA5mf+I
Fcs+gM7EOw6bFA3l1y5tPmRQAhVILRMOyrCtfHI3xv4YOgHN/CEKpBcMgegcAh2U
4IRkWlfqpi6eBN285MqENwb7yfJk/uBMAv3nCgkx43/VC8TrOZSAjl4RYD1dwk2M
B3Df2UcHh26H9/0Y85YgIAf/yk2+EpJvP7BoVAhv2dl+7eUkPcGQIw3+bZqe5DfB
F3xkofLnK9P3uWMDjhn6M6l9GPHK7yW8jgNYrcv3z6qym3ENI9oJ0ejo+n+0NTW9
rGGwyTaXfEUUZ2oHwBvygn9zbgn6aPB0o1dsjGfrO0t+GzsxN8cTqS8SIKuisDpz
vekNBc9ecrctiz52J4jZTZ7y39TyRIn9ZQkPkJL/tI4TSk9V9XKg/+612kT8HIld
zV0NAApwswgMwjkgbGYeAzRCAXzq/3lstIMi1ZXSdxt/ltwbuQBYhK0iIjMgBeT9
OKrFKDkiNOXOPdEYvdcv17DG+bK2NQW5s9IRJEn5rq5H7Pv579LEEMMATQcOTLCk
m4/FlwwVwaGk5Rv3J1sdGK4RcLum+H7McAsUwLWepvUXdgiMX4COs09PpobDcs3i
E0RTVWTLWHhEBKBw+svLypsKoE4xOCpc/ye7qGOxtuN0YtWInklJDAtJReKGJ2MT
4tWWYNmh4w+wkB8nMdBiJJ6NTj6BKYDDYXiousUWhbloawV0ixhI6YTpcmfu+IyU
SKYPcrrvVHu+3LSbuoYz+R0u5QA6VtROl5hEqO5aXhjk1u6xWcJC2d88jeieZarb
zH+8iLkEqvbPfyvZ5NoPrzg85jEj/E7EsNERS464EHycZjyFNT/VxrdPFqWZqj+k
F7yFHTwWSeu4PLV9lHnvPzLwyNAZgcYZuCLi3yDU0f/mVGurcXCWlV9ZT6qq2+Z2
Dv4UPa5f8wcM0paupq9xU3NAN6ngknbS71wNMzUfkhlT8K+plym4gsNJthXagY7R
A8NQqPWYVhNb4ZU6UoFC4usPVSyBpyWv0HDeW/wWCPAnOe7uTUI80a5AnEN+XRJh
mjBiR2fCFumjNASfLpRd3VgI3Yj3pFIxVyzBKe1Auue35r33jKg43f7HfedjDhpY
Ep6c0It+26alvzG4NciLxS5m1MYjA30OTVwWeKGHlaqTsj2CxPExblvhxl5YNXdV
vEQd6BMhPu0yHWlDEgYllZqIuKRvY+xWbnWV/Lyq8dIlnWTQT/oXRvrVXYBXC5Ms
N0DqC65PXRCzJjlWOdKvmfmnTMQhyfq8+3Is2jJ1QcVxBhrUabqb5EDbPqqQOW3M
HYK1cIdUZXJiARIgQ8nJKkd0Ip39EXhhw/zC3Ivxj1RCuDwTSoieWNFjQxD/mhgF
xhlfVRFClM6wzcyix7RJ5LORECuQX+1lWViA937gG+rWCK2JwCkMYIQHJ4vhO+R1
t9Qk8q2YJNA4edw/xu/qaT1/sGKwM0FHy5yV/IREG4IkvkqZsxD3/X6BnztVuath
/WE9Z/zCdaIETY0Cy+u9PdrSzacvNhBR5jtdyr6PWt9YNIPdDLhLUov2+6Z3xxiJ
8uY0ZF2sRDN1R1o0lHXoc+LOHW7eRLEBAsc2RFYgSYYbClTZacPB8nLYNqEoHsjb
/CYop5Rqa3ZuNEEvfnBUcfXHdQZ6sRk0k6QZQbTWCdGGSexHwaCkfdbnLpgTRHfD
EkNiqJjGGBbUHPl/elC1bsgeV0voWSYTvghnXahb9D3j8wfTTaxAtIca1rbzQLXx
HDPqls/GLz/KAXMZWkt/IWv7lijqHuHO3jcfJekcgo3M27pLxZzeJHUQJVMaryWQ
gipMnpjK7i1BL5T4YX9WtvsukaU84EElMrG64LBIXlrvVGa4ar+sfP2/2OQmR7Eh
y4YZJRSNoXP1phhVcsXMLwFtlG3FmAA785jwK2oBsD+FAVGs6ktmds5KZ1Sq3oQP
wmTGgHanhxEGx/odioU1xddq13K3Z7dN+pY1QX8MlLZLgUa2Ya6GDHKPRWs7fYue
0eP6FpNqzEywXm4gIpeY1ZgMNQ5ogXiPOr4kMdyalCLA4FdPggpS2iDApIE11ri4
9OHTUYmMfj+LH7X7R4GYIaZWB8adg9ZPvZpDFywYtLbrnDe4nnRTWRUO9v7eziBo
NeGixTbBdwp22Ra+pRHqNSBHCyqRADYrlTQ9GB9z9c0X2YMtofWzX/rfdgnmIwje
0KAUgiBOb4vYg5aqOXShsWXUhj8ba3S1cejgMq2+5SDcyXB7JQ1YmE03BJOktHql
D8eChBE4KBRs5N2L4x1v6MN7vQrjYQko8amr0xoBrgA5jWU+rfpgMXnDXX9pFIWb
iaHdFzhqtrpfgbNqx2BP1AqI95kaClUiw30GIRwcoxAdMC5MnPNggU6OO8qJ0gJB
mHfx4a9kiCNBMGabLFSjoN0Cb/sL6gmF1Vjx/8ve67PUwO+3z7Bl0pmcXWEt6snQ
lxjBFy8RioIEuc5O6+fG8sJO27a/oQbMi0lI3+hSWV/zlO3FyUZUoz1rxXYE5lXZ
aZOKofHmycqeBiiQz2D17kcOABz5Y01k7SKjibSNgiZVdOfKz10YNf6VILZqqVYH
d7CUzZXEqB3IZm/sujd7fw/WDppfoIHfMOzHYpRlQ7ZCXPerV55wjcKavmhWFb47
q61Kp4H4XhjMn/qQe5JegmPYgt3F/Um8Txom4T9da03zJs7pgjJ5M9T2XP3vq2id
TDBuN65XnyQxOgDDJGX5F15FEjxzDJriWMFjJRDTZLKgLRfQBLmWgp3EOdWwTCU6
3PgCYkuett+Qrl+RyNWhTHX6yTlypUJmt4n0MBMzjXjmgKO7c1D6g9aFev0Zn0BV
my0muLbNZzx827I2dV+O17NJfkZzhM0wu813ebj484biwy+rvSE++mg977KvQWOY
1nqDIrd7KkSUXVb3G9Td257gLxCDPHTizj8tiyVvAkRRNi1/M/Y60ES/RJUYvKin
UXn1HF8cj0fah6KRCzu8P7Ynpb/6Hzy7utoU8ZOBNmhzijjeSJJzrnhdgsKB5WN8
rLKNa8nbPW8dBeW9MZDKRVXVuEVKqrCEg00o+kgM93u4tR3DTCDMI0yTgVQEvNYT
PiS7RUZpeYi1dLshfnVphKKy8mJTsr8raCzhOxdbJipeLbB2HctQMZU1d/x6968S
7yEx4t++7KLqwYBJUpjh2qczVI4bt6S8WzDOQqM/Y0FGJej2nAsmNFatcS6byHFm
B+w/w61aCs1LTW1pQa9rZKbI+UbsfXOFE5OzZuKd9KqjAN8mf4GrJWokE1R5+y76
Ac3rAMo59DdOWoUlZ6W3vBqxIR3v6pbzB2x799VxFNLDLnQEm4veb41BVb56wRSa
8aR7KiaNDvAq+S7ajd9zDsRCLsIUUAtyEIEkGtMbeu6hB4xVJj2CFAewMbqzgLQy
pSLUVPV6+QFk+7YiWs1TRUeABT5MSCdRq/kaqnut+3LzpSAQKY1WwHUE83W19cY8
NR7oA1BUY/efRQdnC9q219yX6klHHgv1tbqpoc4+D127hzcjDRVtzPQQI6Yv5eLP
JdqrKSk/j+iHyvzfdw8kQivYQsIoqlccnwU9nRMZ/5bcbBmKaBs9halEIFVgSpc2
unJ6kYtjX54oJDgXyXKS47KcZYFYWcQbDKTxzr35k6buTzrhAX02nmfb/ntd0jPR
b1GQgFxAyC49Xdfnyb53pSWD/yKtLmWv5Ll6P+Dj7jgWUjXav+3LrPxRaf6pohIS
o4w0FAqJObafItAKhT4x0mzm0ZEfRwv/sgMQw/TbAmJz3Z3gVuQn6geUr9bPacom
l5kvNR3G8ILmgWfKXwozvGEh3UA32GC+JMIHaUTRfMSDF1yop12H2PxHsux+j+3Y
0L71Ky3UR1cyyzTnIQwFGBhYIP62HQpFnDUs1cXAoprQgJ8BSgXDsPwQ2jR6mNW4
vMCE56qtIMHS6N8iDLkjdbxe3xFuFMS09M0HxByLNqZMAgj95POWy/PTdJ9Z0NrX
OglUYvAM2Q1W6YnbJxQzHVk/mpcnb/SrKqoVuytlIwqR4EQ/qdRnAb11uexI6q66
deHValzTUwKDFPcgWywjTFfKvbBekoN4Rbu8siAYTnjR63qoDn+8tgXBXRjtbY4l
JrCF3EYntiNEuP59asJO2CsdX7rmbaGeuVqsJKyEha0Ki/Q1dUb9DkBQN9gBOqWC
vLIsv8XGpoQZtOlYo0iSQ4HEsjg9YAH5yBN2MZYm6aQRKDOw9pvtfCkTfs7ipeDh
HV5J5sYVl2zOCH4OM9VOxWKS2x9fywffer1fYEUTeJmhRnp018WMhHOV/+LnpnMf
kBHB0v+3jkR9IuV5G+nCpVy5v8Dnr45wx9rp9W2/K2o/+KQvvUv+0vVtEZ2KPRtN
18/p/zgWINdKiwcm2IiRWXlFqutOI90+2UTaSxqlFp1s/LXcIU4ALPc+LSRYujaD
C8j19hGm1mfoFQN1A2yd+XY2/MDCvqImzn2P33EAy05YmHNhMeI7UQetHuFJe3gd
4JrxdzaVQye37eskhMAn0negtGc08uX07rmlXU2NmpYsj6TK4Rc+q0kZny1vyWht
oC6YMlhPBY2TkQ6Kw7hkof83RFCBDuGludEkznjKCPGZ802nQlTHRjW+ibDzj+al
WjbD8iUJ+tb2teJvehO9ll3PBwsGaYMugfd+X1dmP16N8TQTuUz0iH803hO+Es/6
HgCpVfXMgRlzDs+015UdSrUpVQsnD+8FS/zoZ9kvEF/vnzf8jPW04ZqGmh4xwekf
6OWKhCn3cUqtQr/mXV1hFUbe4IhYWWvTYmwrTHV//2L6/wOLVr2Qptpy5RiVDaMK
Bp2TeUCe3aCURYMUjh/nT5MFnv+Swn9KHkVyo5E/F+05tkMJltoYAhOTe7UwSpo3
c/y+buA/3/exWOXHjMAk6JVnjyI+0UU4pWoUBmb/PPfR1K/sldEvg3JPXY5D9GcS
whRZP6moqdFcwr2VDygtzJDA6S8n9AbMrrpNkVnDWh+QoMME8SqKxc0UCWpa1TLV
zB1q/JLXuzEM4g1XnrdpXSPNr6lCc42NzCh9cAA6obBqi68Au1XPYRUQAbpFioK0
mhz1UKCNPQ7v539urI2I27wqUfbElkq3QNFf12m4svv93h6MM6MD/Um3fMeWN3ex
pAy/Q5Ne4FQjzSWM3wt6qVXGYJ/jzhLVaf9czZXGMLQvzSamyn9zSvfYxiArVIBY
PGdD099E3O2xieYGtByNOOb0mVniXBQj90LzSCycqd9Xr+N32pK3BJ2Y4WpCbVPw
VADLVXP7QeW/v/SjTiPjdzvJ1woDfw0bHxqGVJSKO4mUSR+/SNx3R/5055V4+mIm
8EHqot4/NXo31mGKLSDfUpFrFdM7lwlxRA4ReZS29vtFW2WdcbRIKx64atua3Tpr
KP4RAiRgK43k5A0Wz0vaVt1N0cZPhdPHSe1DMZo0KdhwG1024Z1ssL3pwgA4QCP+
aMT+Fe6n496om+ylGD0ZbL4YXdMz3kTi+8agzk1PP5oWAWy3Uz399qrbc0G3YMyV
RBOY1tqFzEIuwtge4EWJODJRQd46tCMo4Q69xoy3RCqST+0AcB+n8l5xyOdtv+Yl
5G76L7lX06/uaMVueBal6dRwEQft7mjX8LpYbVOoi27ZkrtM72GCgHSI0DKrRBgl
QuDpRsrXjS+Qh5bqMbP9fTFGyk1GrHP1A2N+HPqsNLpG+1aV+LnLWs2nAzsv99P3
wQbvZyBufuzz6CCtlCx0eXHjqmkruHvNTEnnyevyzUYcGEhkygPyXsW66b3YMYol
sIFwxHbnGI06vxnwoLbuikwB2JBXtCpxoAoRe5pcOexsyf4UHXuSwe42dhLFB2v3
qWyrFzgK4ERPz9o+JW/Lbr4k73e0xiGOhrI3V2BDhGEDF8hVBTTexea/4HZbepJN
CR83r8cWYvAnRp4hWFVgnZXutUvuVAz3i1XD6gG93z2Uc9M7H8icO7BCUaJ2N4n+
ajOMpJ9FEP+rbwqiyT7S06Tyizd6FhhfLjvxXsj3+UQdzOLjDEWVSptagNxaOhaZ
3rKtpSsqkXSgUSb3RiHY7MBRAzU0IQLS05/LfXhBQedDjsVz4PzvkiRdOUSZswix
o7A/5JgbkAPVIVOc+WoLYOFl03/IHT3nyvIVDZnLQjrZbQaHhPCza9ug/bZXmc4p
T7S1LuS6GmsjptE9PX18ymB0J2GgeQ2zFlmtI9hTflF8c6kQ9kJjBX0xxbHxbafd
/bfeqVFrbFPDIgDHxSWWkBE26GKWIgOzAu+bwM4Teecs9j4am4kCXTkNFV4dwFKL
Lg238rSqL4q/hOdEzlFM0SPHeMEx/i+IFwiGGl6BK5x8VVizY2TQ7Ru6olLDUzqR
Lh6yPDIO1B53Ef/4Gom6jpYrJ4nyHWVYbRSA0RnQBpfStoL8IucNhcseA2+w3GLc
driCPTTSUMVEk+TTJkQ55LjhqXsSurOH3hQ6bUKLw4zi1HlzzCWYYGOk7yHjAtgp
QuaW56OuLRs+MrMFKQteD4JVxpZ7KTjDlJOCOtdxtfPMZ6JXkiKXrk+zbKNuSUR7
l4SBwP/slbILIWoTzDcOufr0Tsgl0x6EIojbgm0bENxePTPSVsKN55XpT/rPRgJU
Cw2TYSScMjQFe/K/Bzqn1j1yXnwuQN56DaWFhIT4CY/9ybmOAfaRG780ux1+DESq
uCKb0hPViiLTOyi9jF260c5CeYTVBmmDbK9F9KVCAJHIg1y+hOPQhjjVGa8ebEeK
1G6LjbShPBbWPQJCCggN5ykhQSRinnuym+rS9Xqo6j9N70K+P+LNu5VHJqPMhEZD
r8wxHVE4Zbm9ImOL9Ew7XewRhXCigtNxutOYk9lnaQqPh7Oeehliu/HVWJUt7O97
EDYyZs+vKMxT5UFgcxQ2ztBUEFyZby1yd5i433MrU/by1mWyaEN9SD+5KJ85x7x5
9legCKBs1zuW40QYpiGi5yHoPIRvo8GQADkOXAMxgBSi28+xnGF1iNZf9Ipjh8uo
/lQvw5oNvdK1WirHWBX7zBroFzOge9mHx9yCImOGhTmTpb1OmssaQjFLsByzSAAW
+oE4IAI0D8dXQcLAC9M3YMfFFpCeU+WQbGnmkCyr/14afzo4tVED/pgpeRPnMqly
KIzpn3jPcl+J1aPv1iF7Os8G+W5IfvFi2HxbsG1HcF1j/hEGh4YOqns5Ih2YIeja
BXUYkeczHzCLuVPA1/4zvZx7NwsvbbvhXZUa/BXrZk9L0vbox9gKO3BuLD+p+Pxf
jOXEq4XzoEff9Mqrp5xWWmD+nblkKAsZQAqJUKThxjqB4c4GZZuOHR0f8Xp4MhFQ
60ctkL7u6ZP6/GWF61zZ0RcqUvXlYXD7t1kB/mBvczIg0AOKR/xKZBVgnFbP6p09
4ysmXNazHYS4z85xVg5jo8Tlmu+rLVv+mjf/M1AlRiax63rmOnKdVZ4dqIveig2B
sqzsH7muwqgjuJX9ZfO5zdvsMDnTYErzOXB3osaRbnAc5ND8BCoNAQ4YwjwQNz7t
SuUR66z33JB8mh/OY0DLP/bi5HJeDmfsmaumCP93QXp+YwTeeVeC/7uBQSnPwymv
0u0L5geZ1f4FRz09EvGJbzQiHzfQTNNWDOCjUb3XQHvY86LnTLmeXFZeMJQGDe/i
TQFn5a6qS88nzdxHTqbiEL3VBXKGQf6dh4B4blOiiAbPNEihdtrXSh200CqqEOLm
o0oc8mJfe2mtFOswiLrfuy8ARF+gTBmu3eZDMSDqe8gcuXiHvHVTNabzlinriTsY
Du7bmULCG6E+8QNfBZnrIG9i/YFmnYcpyQsnm4rrEtEOBSsX1Z3fjOWDVqX/ZAED
m0sf2XV07181qpUBfl1jDpfwlIhyvh4MOjIKRWYdR+bKJ/bNY6/gWkQa/gLIl0GH
sj18DxNeFtDAbHa/z84lV4Y0grJmaOSVB4o8pw2o0Yxeir1CYoLMXLDDJNI+JZQ/
LaHyv+7tRSgElmcr25IeZlJsWXSXivluZ97Tnwp1aO4gh/IoYrVz7SlLly4M8f0p
2sWObWhNtFWiwsWKMl0Tf4Ou6seJFqqnMXNuhJ3fjCyeMD8to2NbhBL8/muWxztw
Y2Jx3c7XHZGTm67M1CtbIr5X4Ojh5BjqnNVyeTlkjajeDlzraD147GWyPf5AhUtm
1yN9cIv45KsjpoQg1VQNQ6WQ7ZrsGEltEt/ahYvWkvH44mnVCziwGFDa0bBNCa7P
gMrq1kzoa1T3FCFtdjwCuMnEBgYaqsyYoLaQzawA6WsTAWVdbRI7EHm+yc42dcmE
upHc/ZTV1k0oOC+MEkXscRC/UHMOVNSWEZ5YQRgzWAGV33PNH6voveI6+x6XcMvF
W1Dr/9YjaK4vL/5Fl4OvxDkoLlWGkt/g7DX5a3zNYzG9puGvou0OCBTnYIg7EBIO
GI04eq/0ZgrGOcr0U+skV7MMbHBhFhNxs+YzTrWY6G/Uz61Dsh+64aOONlVlY7ly
fopvUk/XfZBO6OZuWOri5w8SwaD4mkti9BvDfo2QmmIDRVnMtRozmPZ31St4u2jx
/J3VuJU/RqsH/bxNqPuu2HZRqBfaF6CkQznFaETXc8Kl8+g1kebl9cLUhGESUDqK
qwd6eAUC0bSx/qiLh1KMwLjbVwqvlze42XD98F9FZfbIiMYjhxaJNdhYk+d+ra/f
vhFfgs+FrSYQfRFILmTylYzZBtBOK8kMQFXyYyn3ZKRT6euWrgi05xu97fjQa7dw
4xgggmydkmF81VJLx92/T9EnEtkxH7oVafU6TqbO+Y9YNBaxWwIv5efmGXwTcOI2
o8MLMnWn6i45bQUMHGX80nidqg0DK986amtYGgXfXVjKKokbDLU+55zuHjd6NNgj
Ga8FYSjdYeNldctuVacDEKstR/7dgmZBEVwvzxjS4zsnc2fiXzPCJww9vTm1C6Kp
p4yA6JQwPwpC+y3+LcaCo81tyQpOsEYxFdEIxt2m48Mc07VID5LpqS5ZVsd8D1e1
oNBvamBm1mCuSgCD7d6+xHFOzKuMTpSc54Y6Jv3l/YdxRgzlPSsz3jOhQc3HitLn
4+ncl11kBABG4EWy/djQqo/BekJ0tEFeOLxX9i8NaCEsObRGbitZX8pN/qdxQ75p
UBXBOMUeC1lv6OV5waTOfTRGp8S+PsCPMq/YQS0Uad4V3kkInzrYhynnpElmsil5
tr7RGhrejjDCOeqB7GhuPLw6WfhAF+DoDIa0kGrSxOGjEuFt+kGH3AUfGyRWbuUz
yLgEVC+5epTKcogKUn8PGIY5s0Ra8wQggKXQwr241ErannZ3C2/mT+1UXSYoJJ7c
lWrktWxXV6pGyO5Ri6HqxyDMEHZUhuDcbcHo1Aoo4Bl6e+kEEdryqo7RyVd8xKsy
L5oaksAyfsFxzqiq1FvSrMudpI85jyKcjP3FBrcIntYTWdm9GT+0s6ZwUJQ54FFC
CvfUhHEQjLojEu+7GOCN9kPYgctaEQP0zh3qiGRvilRRDNvqTgoZqsBUQyuecKHc
n3ts1e1VvInqkneIlA1akBdaD47KLPo1c4JMVg8mdMFCOjISP1NDEIMFVPVZwMuc
VhabfuMA4s36Xl6lJtCO1J+aFasTh/qgCeLQGEKEsjA4/7imbPkvXHCYk2eP55T1
gjEXsgJy1lrSS9AEiskhwUeKCfSIlfY5p/iMW5pZbEXPIk8VjsP8QJg9F/6qVJEu
cFRl6y79yMsoJITE/zPtXfvvlNP2PTzcfHX6U78tF6g=
`protect END_PROTECTED
